magic
tech sky130A
magscale 1 2
timestamp 1647745527
<< checkpaint >>
rect -1266 2308 2814 9166
rect -1266 -1091 1554 2308
<< nwell >>
rect 294 3632 1254 7906
<< pwell >>
rect 378 3201 654 3589
rect 894 3201 1170 3589
rect 378 1975 654 2363
rect 894 1975 1170 2363
rect 378 1501 654 1889
rect 894 1501 1170 1889
rect 356 169 1192 621
<< nmos >>
rect 458 3227 488 3563
rect 544 3227 574 3563
rect 974 3227 1004 3563
rect 1060 3227 1090 3563
rect 458 2001 488 2337
rect 544 2001 574 2337
rect 974 2001 1004 2337
rect 1060 2001 1090 2337
rect 458 1527 488 1863
rect 544 1527 574 1863
rect 974 1527 1004 1863
rect 1060 1527 1090 1863
<< pmos >>
rect 458 6503 488 6703
rect 544 6503 574 6703
rect 974 6503 1004 6703
rect 1060 6503 1090 6703
rect 458 5061 488 5261
rect 544 5061 574 5261
rect 974 5061 1004 5261
rect 1060 5061 1090 5261
rect 458 3701 488 4101
rect 544 3701 574 4101
rect 974 3701 1004 4101
rect 1060 3701 1090 4101
<< ndiff >>
rect 404 3548 458 3563
rect 404 3514 413 3548
rect 447 3514 458 3548
rect 404 3480 458 3514
rect 404 3446 413 3480
rect 447 3446 458 3480
rect 404 3412 458 3446
rect 404 3378 413 3412
rect 447 3378 458 3412
rect 404 3344 458 3378
rect 404 3310 413 3344
rect 447 3310 458 3344
rect 404 3276 458 3310
rect 404 3242 413 3276
rect 447 3242 458 3276
rect 404 3227 458 3242
rect 488 3548 544 3563
rect 488 3514 499 3548
rect 533 3514 544 3548
rect 488 3480 544 3514
rect 488 3446 499 3480
rect 533 3446 544 3480
rect 488 3412 544 3446
rect 488 3378 499 3412
rect 533 3378 544 3412
rect 488 3344 544 3378
rect 488 3310 499 3344
rect 533 3310 544 3344
rect 488 3276 544 3310
rect 488 3242 499 3276
rect 533 3242 544 3276
rect 488 3227 544 3242
rect 574 3548 628 3563
rect 574 3514 585 3548
rect 619 3514 628 3548
rect 574 3480 628 3514
rect 574 3446 585 3480
rect 619 3446 628 3480
rect 574 3412 628 3446
rect 574 3378 585 3412
rect 619 3378 628 3412
rect 574 3344 628 3378
rect 574 3310 585 3344
rect 619 3310 628 3344
rect 574 3276 628 3310
rect 574 3242 585 3276
rect 619 3242 628 3276
rect 574 3227 628 3242
rect 920 3548 974 3563
rect 920 3514 929 3548
rect 963 3514 974 3548
rect 920 3480 974 3514
rect 920 3446 929 3480
rect 963 3446 974 3480
rect 920 3412 974 3446
rect 920 3378 929 3412
rect 963 3378 974 3412
rect 920 3344 974 3378
rect 920 3310 929 3344
rect 963 3310 974 3344
rect 920 3276 974 3310
rect 920 3242 929 3276
rect 963 3242 974 3276
rect 920 3227 974 3242
rect 1004 3548 1060 3563
rect 1004 3514 1015 3548
rect 1049 3514 1060 3548
rect 1004 3480 1060 3514
rect 1004 3446 1015 3480
rect 1049 3446 1060 3480
rect 1004 3412 1060 3446
rect 1004 3378 1015 3412
rect 1049 3378 1060 3412
rect 1004 3344 1060 3378
rect 1004 3310 1015 3344
rect 1049 3310 1060 3344
rect 1004 3276 1060 3310
rect 1004 3242 1015 3276
rect 1049 3242 1060 3276
rect 1004 3227 1060 3242
rect 1090 3548 1144 3563
rect 1090 3514 1101 3548
rect 1135 3514 1144 3548
rect 1090 3480 1144 3514
rect 1090 3446 1101 3480
rect 1135 3446 1144 3480
rect 1090 3412 1144 3446
rect 1090 3378 1101 3412
rect 1135 3378 1144 3412
rect 1090 3344 1144 3378
rect 1090 3310 1101 3344
rect 1135 3310 1144 3344
rect 1090 3276 1144 3310
rect 1090 3242 1101 3276
rect 1135 3242 1144 3276
rect 1090 3227 1144 3242
rect 404 2322 458 2337
rect 404 2288 413 2322
rect 447 2288 458 2322
rect 404 2254 458 2288
rect 404 2220 413 2254
rect 447 2220 458 2254
rect 404 2186 458 2220
rect 404 2152 413 2186
rect 447 2152 458 2186
rect 404 2118 458 2152
rect 404 2084 413 2118
rect 447 2084 458 2118
rect 404 2050 458 2084
rect 404 2016 413 2050
rect 447 2016 458 2050
rect 404 2001 458 2016
rect 488 2322 544 2337
rect 488 2288 499 2322
rect 533 2288 544 2322
rect 488 2254 544 2288
rect 488 2220 499 2254
rect 533 2220 544 2254
rect 488 2186 544 2220
rect 488 2152 499 2186
rect 533 2152 544 2186
rect 488 2118 544 2152
rect 488 2084 499 2118
rect 533 2084 544 2118
rect 488 2050 544 2084
rect 488 2016 499 2050
rect 533 2016 544 2050
rect 488 2001 544 2016
rect 574 2322 628 2337
rect 574 2288 585 2322
rect 619 2288 628 2322
rect 574 2254 628 2288
rect 574 2220 585 2254
rect 619 2220 628 2254
rect 574 2186 628 2220
rect 574 2152 585 2186
rect 619 2152 628 2186
rect 574 2118 628 2152
rect 574 2084 585 2118
rect 619 2084 628 2118
rect 574 2050 628 2084
rect 574 2016 585 2050
rect 619 2016 628 2050
rect 574 2001 628 2016
rect 920 2322 974 2337
rect 920 2288 929 2322
rect 963 2288 974 2322
rect 920 2254 974 2288
rect 920 2220 929 2254
rect 963 2220 974 2254
rect 920 2186 974 2220
rect 920 2152 929 2186
rect 963 2152 974 2186
rect 920 2118 974 2152
rect 920 2084 929 2118
rect 963 2084 974 2118
rect 920 2050 974 2084
rect 920 2016 929 2050
rect 963 2016 974 2050
rect 920 2001 974 2016
rect 1004 2322 1060 2337
rect 1004 2288 1015 2322
rect 1049 2288 1060 2322
rect 1004 2254 1060 2288
rect 1004 2220 1015 2254
rect 1049 2220 1060 2254
rect 1004 2186 1060 2220
rect 1004 2152 1015 2186
rect 1049 2152 1060 2186
rect 1004 2118 1060 2152
rect 1004 2084 1015 2118
rect 1049 2084 1060 2118
rect 1004 2050 1060 2084
rect 1004 2016 1015 2050
rect 1049 2016 1060 2050
rect 1004 2001 1060 2016
rect 1090 2322 1144 2337
rect 1090 2288 1101 2322
rect 1135 2288 1144 2322
rect 1090 2254 1144 2288
rect 1090 2220 1101 2254
rect 1135 2220 1144 2254
rect 1090 2186 1144 2220
rect 1090 2152 1101 2186
rect 1135 2152 1144 2186
rect 1090 2118 1144 2152
rect 1090 2084 1101 2118
rect 1135 2084 1144 2118
rect 1090 2050 1144 2084
rect 1090 2016 1101 2050
rect 1135 2016 1144 2050
rect 1090 2001 1144 2016
rect 404 1848 458 1863
rect 404 1814 413 1848
rect 447 1814 458 1848
rect 404 1780 458 1814
rect 404 1746 413 1780
rect 447 1746 458 1780
rect 404 1712 458 1746
rect 404 1678 413 1712
rect 447 1678 458 1712
rect 404 1644 458 1678
rect 404 1610 413 1644
rect 447 1610 458 1644
rect 404 1576 458 1610
rect 404 1542 413 1576
rect 447 1542 458 1576
rect 404 1527 458 1542
rect 488 1848 544 1863
rect 488 1814 499 1848
rect 533 1814 544 1848
rect 488 1780 544 1814
rect 488 1746 499 1780
rect 533 1746 544 1780
rect 488 1712 544 1746
rect 488 1678 499 1712
rect 533 1678 544 1712
rect 488 1644 544 1678
rect 488 1610 499 1644
rect 533 1610 544 1644
rect 488 1576 544 1610
rect 488 1542 499 1576
rect 533 1542 544 1576
rect 488 1527 544 1542
rect 574 1848 628 1863
rect 574 1814 585 1848
rect 619 1814 628 1848
rect 574 1780 628 1814
rect 574 1746 585 1780
rect 619 1746 628 1780
rect 574 1712 628 1746
rect 574 1678 585 1712
rect 619 1678 628 1712
rect 574 1644 628 1678
rect 574 1610 585 1644
rect 619 1610 628 1644
rect 574 1576 628 1610
rect 574 1542 585 1576
rect 619 1542 628 1576
rect 574 1527 628 1542
rect 920 1848 974 1863
rect 920 1814 929 1848
rect 963 1814 974 1848
rect 920 1780 974 1814
rect 920 1746 929 1780
rect 963 1746 974 1780
rect 920 1712 974 1746
rect 920 1678 929 1712
rect 963 1678 974 1712
rect 920 1644 974 1678
rect 920 1610 929 1644
rect 963 1610 974 1644
rect 920 1576 974 1610
rect 920 1542 929 1576
rect 963 1542 974 1576
rect 920 1527 974 1542
rect 1004 1848 1060 1863
rect 1004 1814 1015 1848
rect 1049 1814 1060 1848
rect 1004 1780 1060 1814
rect 1004 1746 1015 1780
rect 1049 1746 1060 1780
rect 1004 1712 1060 1746
rect 1004 1678 1015 1712
rect 1049 1678 1060 1712
rect 1004 1644 1060 1678
rect 1004 1610 1015 1644
rect 1049 1610 1060 1644
rect 1004 1576 1060 1610
rect 1004 1542 1015 1576
rect 1049 1542 1060 1576
rect 1004 1527 1060 1542
rect 1090 1848 1144 1863
rect 1090 1814 1101 1848
rect 1135 1814 1144 1848
rect 1090 1780 1144 1814
rect 1090 1746 1101 1780
rect 1135 1746 1144 1780
rect 1090 1712 1144 1746
rect 1090 1678 1101 1712
rect 1135 1678 1144 1712
rect 1090 1644 1144 1678
rect 1090 1610 1101 1644
rect 1135 1610 1144 1644
rect 1090 1576 1144 1610
rect 1090 1542 1101 1576
rect 1135 1542 1144 1576
rect 1090 1527 1144 1542
<< pdiff >>
rect 404 6688 458 6703
rect 404 6654 413 6688
rect 447 6654 458 6688
rect 404 6620 458 6654
rect 404 6586 413 6620
rect 447 6586 458 6620
rect 404 6552 458 6586
rect 404 6518 413 6552
rect 447 6518 458 6552
rect 404 6503 458 6518
rect 488 6688 544 6703
rect 488 6654 499 6688
rect 533 6654 544 6688
rect 488 6620 544 6654
rect 488 6586 499 6620
rect 533 6586 544 6620
rect 488 6552 544 6586
rect 488 6518 499 6552
rect 533 6518 544 6552
rect 488 6503 544 6518
rect 574 6688 628 6703
rect 574 6654 585 6688
rect 619 6654 628 6688
rect 574 6620 628 6654
rect 574 6586 585 6620
rect 619 6586 628 6620
rect 574 6552 628 6586
rect 574 6518 585 6552
rect 619 6518 628 6552
rect 574 6503 628 6518
rect 920 6688 974 6703
rect 920 6654 929 6688
rect 963 6654 974 6688
rect 920 6620 974 6654
rect 920 6586 929 6620
rect 963 6586 974 6620
rect 920 6552 974 6586
rect 920 6518 929 6552
rect 963 6518 974 6552
rect 920 6503 974 6518
rect 1004 6688 1060 6703
rect 1004 6654 1015 6688
rect 1049 6654 1060 6688
rect 1004 6620 1060 6654
rect 1004 6586 1015 6620
rect 1049 6586 1060 6620
rect 1004 6552 1060 6586
rect 1004 6518 1015 6552
rect 1049 6518 1060 6552
rect 1004 6503 1060 6518
rect 1090 6688 1144 6703
rect 1090 6654 1101 6688
rect 1135 6654 1144 6688
rect 1090 6620 1144 6654
rect 1090 6586 1101 6620
rect 1135 6586 1144 6620
rect 1090 6552 1144 6586
rect 1090 6518 1101 6552
rect 1135 6518 1144 6552
rect 1090 6503 1144 6518
rect 404 5246 458 5261
rect 404 5212 413 5246
rect 447 5212 458 5246
rect 404 5178 458 5212
rect 404 5144 413 5178
rect 447 5144 458 5178
rect 404 5110 458 5144
rect 404 5076 413 5110
rect 447 5076 458 5110
rect 404 5061 458 5076
rect 488 5246 544 5261
rect 488 5212 499 5246
rect 533 5212 544 5246
rect 488 5178 544 5212
rect 488 5144 499 5178
rect 533 5144 544 5178
rect 488 5110 544 5144
rect 488 5076 499 5110
rect 533 5076 544 5110
rect 488 5061 544 5076
rect 574 5246 628 5261
rect 574 5212 585 5246
rect 619 5212 628 5246
rect 574 5178 628 5212
rect 574 5144 585 5178
rect 619 5144 628 5178
rect 574 5110 628 5144
rect 574 5076 585 5110
rect 619 5076 628 5110
rect 574 5061 628 5076
rect 920 5246 974 5261
rect 920 5212 929 5246
rect 963 5212 974 5246
rect 920 5178 974 5212
rect 920 5144 929 5178
rect 963 5144 974 5178
rect 920 5110 974 5144
rect 920 5076 929 5110
rect 963 5076 974 5110
rect 920 5061 974 5076
rect 1004 5246 1060 5261
rect 1004 5212 1015 5246
rect 1049 5212 1060 5246
rect 1004 5178 1060 5212
rect 1004 5144 1015 5178
rect 1049 5144 1060 5178
rect 1004 5110 1060 5144
rect 1004 5076 1015 5110
rect 1049 5076 1060 5110
rect 1004 5061 1060 5076
rect 1090 5246 1144 5261
rect 1090 5212 1101 5246
rect 1135 5212 1144 5246
rect 1090 5178 1144 5212
rect 1090 5144 1101 5178
rect 1135 5144 1144 5178
rect 1090 5110 1144 5144
rect 1090 5076 1101 5110
rect 1135 5076 1144 5110
rect 1090 5061 1144 5076
rect 404 4088 458 4101
rect 404 4054 413 4088
rect 447 4054 458 4088
rect 404 4020 458 4054
rect 404 3986 413 4020
rect 447 3986 458 4020
rect 404 3952 458 3986
rect 404 3918 413 3952
rect 447 3918 458 3952
rect 404 3884 458 3918
rect 404 3850 413 3884
rect 447 3850 458 3884
rect 404 3816 458 3850
rect 404 3782 413 3816
rect 447 3782 458 3816
rect 404 3748 458 3782
rect 404 3714 413 3748
rect 447 3714 458 3748
rect 404 3701 458 3714
rect 488 4088 544 4101
rect 488 4054 499 4088
rect 533 4054 544 4088
rect 488 4020 544 4054
rect 488 3986 499 4020
rect 533 3986 544 4020
rect 488 3952 544 3986
rect 488 3918 499 3952
rect 533 3918 544 3952
rect 488 3884 544 3918
rect 488 3850 499 3884
rect 533 3850 544 3884
rect 488 3816 544 3850
rect 488 3782 499 3816
rect 533 3782 544 3816
rect 488 3748 544 3782
rect 488 3714 499 3748
rect 533 3714 544 3748
rect 488 3701 544 3714
rect 574 4088 628 4101
rect 574 4054 585 4088
rect 619 4054 628 4088
rect 574 4020 628 4054
rect 574 3986 585 4020
rect 619 3986 628 4020
rect 574 3952 628 3986
rect 574 3918 585 3952
rect 619 3918 628 3952
rect 574 3884 628 3918
rect 574 3850 585 3884
rect 619 3850 628 3884
rect 574 3816 628 3850
rect 574 3782 585 3816
rect 619 3782 628 3816
rect 574 3748 628 3782
rect 574 3714 585 3748
rect 619 3714 628 3748
rect 574 3701 628 3714
rect 920 4088 974 4101
rect 920 4054 929 4088
rect 963 4054 974 4088
rect 920 4020 974 4054
rect 920 3986 929 4020
rect 963 3986 974 4020
rect 920 3952 974 3986
rect 920 3918 929 3952
rect 963 3918 974 3952
rect 920 3884 974 3918
rect 920 3850 929 3884
rect 963 3850 974 3884
rect 920 3816 974 3850
rect 920 3782 929 3816
rect 963 3782 974 3816
rect 920 3748 974 3782
rect 920 3714 929 3748
rect 963 3714 974 3748
rect 920 3701 974 3714
rect 1004 4088 1060 4101
rect 1004 4054 1015 4088
rect 1049 4054 1060 4088
rect 1004 4020 1060 4054
rect 1004 3986 1015 4020
rect 1049 3986 1060 4020
rect 1004 3952 1060 3986
rect 1004 3918 1015 3952
rect 1049 3918 1060 3952
rect 1004 3884 1060 3918
rect 1004 3850 1015 3884
rect 1049 3850 1060 3884
rect 1004 3816 1060 3850
rect 1004 3782 1015 3816
rect 1049 3782 1060 3816
rect 1004 3748 1060 3782
rect 1004 3714 1015 3748
rect 1049 3714 1060 3748
rect 1004 3701 1060 3714
rect 1090 4088 1144 4101
rect 1090 4054 1101 4088
rect 1135 4054 1144 4088
rect 1090 4020 1144 4054
rect 1090 3986 1101 4020
rect 1135 3986 1144 4020
rect 1090 3952 1144 3986
rect 1090 3918 1101 3952
rect 1135 3918 1144 3952
rect 1090 3884 1144 3918
rect 1090 3850 1101 3884
rect 1135 3850 1144 3884
rect 1090 3816 1144 3850
rect 1090 3782 1101 3816
rect 1135 3782 1144 3816
rect 1090 3748 1144 3782
rect 1090 3714 1101 3748
rect 1135 3714 1144 3748
rect 1090 3701 1144 3714
<< ndiffc >>
rect 413 3514 447 3548
rect 413 3446 447 3480
rect 413 3378 447 3412
rect 413 3310 447 3344
rect 413 3242 447 3276
rect 499 3514 533 3548
rect 499 3446 533 3480
rect 499 3378 533 3412
rect 499 3310 533 3344
rect 499 3242 533 3276
rect 585 3514 619 3548
rect 585 3446 619 3480
rect 585 3378 619 3412
rect 585 3310 619 3344
rect 585 3242 619 3276
rect 929 3514 963 3548
rect 929 3446 963 3480
rect 929 3378 963 3412
rect 929 3310 963 3344
rect 929 3242 963 3276
rect 1015 3514 1049 3548
rect 1015 3446 1049 3480
rect 1015 3378 1049 3412
rect 1015 3310 1049 3344
rect 1015 3242 1049 3276
rect 1101 3514 1135 3548
rect 1101 3446 1135 3480
rect 1101 3378 1135 3412
rect 1101 3310 1135 3344
rect 1101 3242 1135 3276
rect 413 2288 447 2322
rect 413 2220 447 2254
rect 413 2152 447 2186
rect 413 2084 447 2118
rect 413 2016 447 2050
rect 499 2288 533 2322
rect 499 2220 533 2254
rect 499 2152 533 2186
rect 499 2084 533 2118
rect 499 2016 533 2050
rect 585 2288 619 2322
rect 585 2220 619 2254
rect 585 2152 619 2186
rect 585 2084 619 2118
rect 585 2016 619 2050
rect 929 2288 963 2322
rect 929 2220 963 2254
rect 929 2152 963 2186
rect 929 2084 963 2118
rect 929 2016 963 2050
rect 1015 2288 1049 2322
rect 1015 2220 1049 2254
rect 1015 2152 1049 2186
rect 1015 2084 1049 2118
rect 1015 2016 1049 2050
rect 1101 2288 1135 2322
rect 1101 2220 1135 2254
rect 1101 2152 1135 2186
rect 1101 2084 1135 2118
rect 1101 2016 1135 2050
rect 413 1814 447 1848
rect 413 1746 447 1780
rect 413 1678 447 1712
rect 413 1610 447 1644
rect 413 1542 447 1576
rect 499 1814 533 1848
rect 499 1746 533 1780
rect 499 1678 533 1712
rect 499 1610 533 1644
rect 499 1542 533 1576
rect 585 1814 619 1848
rect 585 1746 619 1780
rect 585 1678 619 1712
rect 585 1610 619 1644
rect 585 1542 619 1576
rect 929 1814 963 1848
rect 929 1746 963 1780
rect 929 1678 963 1712
rect 929 1610 963 1644
rect 929 1542 963 1576
rect 1015 1814 1049 1848
rect 1015 1746 1049 1780
rect 1015 1678 1049 1712
rect 1015 1610 1049 1644
rect 1015 1542 1049 1576
rect 1101 1814 1135 1848
rect 1101 1746 1135 1780
rect 1101 1678 1135 1712
rect 1101 1610 1135 1644
rect 1101 1542 1135 1576
<< pdiffc >>
rect 413 6654 447 6688
rect 413 6586 447 6620
rect 413 6518 447 6552
rect 499 6654 533 6688
rect 499 6586 533 6620
rect 499 6518 533 6552
rect 585 6654 619 6688
rect 585 6586 619 6620
rect 585 6518 619 6552
rect 929 6654 963 6688
rect 929 6586 963 6620
rect 929 6518 963 6552
rect 1015 6654 1049 6688
rect 1015 6586 1049 6620
rect 1015 6518 1049 6552
rect 1101 6654 1135 6688
rect 1101 6586 1135 6620
rect 1101 6518 1135 6552
rect 413 5212 447 5246
rect 413 5144 447 5178
rect 413 5076 447 5110
rect 499 5212 533 5246
rect 499 5144 533 5178
rect 499 5076 533 5110
rect 585 5212 619 5246
rect 585 5144 619 5178
rect 585 5076 619 5110
rect 929 5212 963 5246
rect 929 5144 963 5178
rect 929 5076 963 5110
rect 1015 5212 1049 5246
rect 1015 5144 1049 5178
rect 1015 5076 1049 5110
rect 1101 5212 1135 5246
rect 1101 5144 1135 5178
rect 1101 5076 1135 5110
rect 413 4054 447 4088
rect 413 3986 447 4020
rect 413 3918 447 3952
rect 413 3850 447 3884
rect 413 3782 447 3816
rect 413 3714 447 3748
rect 499 4054 533 4088
rect 499 3986 533 4020
rect 499 3918 533 3952
rect 499 3850 533 3884
rect 499 3782 533 3816
rect 499 3714 533 3748
rect 585 4054 619 4088
rect 585 3986 619 4020
rect 585 3918 619 3952
rect 585 3850 619 3884
rect 585 3782 619 3816
rect 585 3714 619 3748
rect 929 4054 963 4088
rect 929 3986 963 4020
rect 929 3918 963 3952
rect 929 3850 963 3884
rect 929 3782 963 3816
rect 929 3714 963 3748
rect 1015 4054 1049 4088
rect 1015 3986 1049 4020
rect 1015 3918 1049 3952
rect 1015 3850 1049 3884
rect 1015 3782 1049 3816
rect 1015 3714 1049 3748
rect 1101 4054 1135 4088
rect 1101 3986 1135 4020
rect 1101 3918 1135 3952
rect 1101 3850 1135 3884
rect 1101 3782 1135 3816
rect 1101 3714 1135 3748
<< psubdiff >>
rect 382 582 1166 595
rect 382 548 413 582
rect 447 548 499 582
rect 533 548 585 582
rect 619 548 671 582
rect 705 548 757 582
rect 791 548 843 582
rect 877 548 929 582
rect 963 548 1015 582
rect 1049 548 1101 582
rect 1135 548 1166 582
rect 382 514 1166 548
rect 382 480 413 514
rect 447 480 499 514
rect 533 480 585 514
rect 619 480 671 514
rect 705 480 757 514
rect 791 480 843 514
rect 877 480 929 514
rect 963 480 1015 514
rect 1049 480 1101 514
rect 1135 480 1166 514
rect 382 446 1166 480
rect 382 412 413 446
rect 447 412 499 446
rect 533 412 585 446
rect 619 412 671 446
rect 705 412 757 446
rect 791 412 843 446
rect 877 412 929 446
rect 963 412 1015 446
rect 1049 412 1101 446
rect 1135 412 1166 446
rect 382 378 1166 412
rect 382 344 413 378
rect 447 344 499 378
rect 533 344 585 378
rect 619 344 671 378
rect 705 344 757 378
rect 791 344 843 378
rect 877 344 929 378
rect 963 344 1015 378
rect 1049 344 1101 378
rect 1135 344 1166 378
rect 382 310 1166 344
rect 382 276 413 310
rect 447 276 499 310
rect 533 276 585 310
rect 619 276 671 310
rect 705 276 757 310
rect 791 276 843 310
rect 877 276 929 310
rect 963 276 1015 310
rect 1049 276 1101 310
rect 1135 276 1166 310
rect 382 242 1166 276
rect 382 208 413 242
rect 447 208 499 242
rect 533 208 585 242
rect 619 208 671 242
rect 705 208 757 242
rect 791 208 843 242
rect 877 208 929 242
rect 963 208 1015 242
rect 1049 208 1101 242
rect 1135 208 1166 242
rect 382 195 1166 208
<< nsubdiff >>
rect 382 7698 1166 7713
rect 382 7664 413 7698
rect 447 7664 499 7698
rect 533 7664 585 7698
rect 619 7664 671 7698
rect 705 7664 757 7698
rect 791 7664 843 7698
rect 877 7664 929 7698
rect 963 7664 1015 7698
rect 1049 7664 1101 7698
rect 1135 7664 1166 7698
rect 382 7630 1166 7664
rect 382 7596 413 7630
rect 447 7596 499 7630
rect 533 7596 585 7630
rect 619 7596 671 7630
rect 705 7596 757 7630
rect 791 7596 843 7630
rect 877 7596 929 7630
rect 963 7596 1015 7630
rect 1049 7596 1101 7630
rect 1135 7596 1166 7630
rect 382 7562 1166 7596
rect 382 7528 413 7562
rect 447 7528 499 7562
rect 533 7528 585 7562
rect 619 7528 671 7562
rect 705 7528 757 7562
rect 791 7528 843 7562
rect 877 7528 929 7562
rect 963 7528 1015 7562
rect 1049 7528 1101 7562
rect 1135 7528 1166 7562
rect 382 7494 1166 7528
rect 382 7460 413 7494
rect 447 7460 499 7494
rect 533 7460 585 7494
rect 619 7460 671 7494
rect 705 7460 757 7494
rect 791 7460 843 7494
rect 877 7460 929 7494
rect 963 7460 1015 7494
rect 1049 7460 1101 7494
rect 1135 7460 1166 7494
rect 382 7426 1166 7460
rect 382 7392 413 7426
rect 447 7392 499 7426
rect 533 7392 585 7426
rect 619 7392 671 7426
rect 705 7392 757 7426
rect 791 7392 843 7426
rect 877 7392 929 7426
rect 963 7392 1015 7426
rect 1049 7392 1101 7426
rect 1135 7392 1166 7426
rect 382 7377 1166 7392
<< psubdiffcont >>
rect 413 548 447 582
rect 499 548 533 582
rect 585 548 619 582
rect 671 548 705 582
rect 757 548 791 582
rect 843 548 877 582
rect 929 548 963 582
rect 1015 548 1049 582
rect 1101 548 1135 582
rect 413 480 447 514
rect 499 480 533 514
rect 585 480 619 514
rect 671 480 705 514
rect 757 480 791 514
rect 843 480 877 514
rect 929 480 963 514
rect 1015 480 1049 514
rect 1101 480 1135 514
rect 413 412 447 446
rect 499 412 533 446
rect 585 412 619 446
rect 671 412 705 446
rect 757 412 791 446
rect 843 412 877 446
rect 929 412 963 446
rect 1015 412 1049 446
rect 1101 412 1135 446
rect 413 344 447 378
rect 499 344 533 378
rect 585 344 619 378
rect 671 344 705 378
rect 757 344 791 378
rect 843 344 877 378
rect 929 344 963 378
rect 1015 344 1049 378
rect 1101 344 1135 378
rect 413 276 447 310
rect 499 276 533 310
rect 585 276 619 310
rect 671 276 705 310
rect 757 276 791 310
rect 843 276 877 310
rect 929 276 963 310
rect 1015 276 1049 310
rect 1101 276 1135 310
rect 413 208 447 242
rect 499 208 533 242
rect 585 208 619 242
rect 671 208 705 242
rect 757 208 791 242
rect 843 208 877 242
rect 929 208 963 242
rect 1015 208 1049 242
rect 1101 208 1135 242
<< nsubdiffcont >>
rect 413 7664 447 7698
rect 499 7664 533 7698
rect 585 7664 619 7698
rect 671 7664 705 7698
rect 757 7664 791 7698
rect 843 7664 877 7698
rect 929 7664 963 7698
rect 1015 7664 1049 7698
rect 1101 7664 1135 7698
rect 413 7596 447 7630
rect 499 7596 533 7630
rect 585 7596 619 7630
rect 671 7596 705 7630
rect 757 7596 791 7630
rect 843 7596 877 7630
rect 929 7596 963 7630
rect 1015 7596 1049 7630
rect 1101 7596 1135 7630
rect 413 7528 447 7562
rect 499 7528 533 7562
rect 585 7528 619 7562
rect 671 7528 705 7562
rect 757 7528 791 7562
rect 843 7528 877 7562
rect 929 7528 963 7562
rect 1015 7528 1049 7562
rect 1101 7528 1135 7562
rect 413 7460 447 7494
rect 499 7460 533 7494
rect 585 7460 619 7494
rect 671 7460 705 7494
rect 757 7460 791 7494
rect 843 7460 877 7494
rect 929 7460 963 7494
rect 1015 7460 1049 7494
rect 1101 7460 1135 7494
rect 413 7392 447 7426
rect 499 7392 533 7426
rect 585 7392 619 7426
rect 671 7392 705 7426
rect 757 7392 791 7426
rect 843 7392 877 7426
rect 929 7392 963 7426
rect 1015 7392 1049 7426
rect 1101 7392 1135 7426
<< poly >>
rect 458 6703 488 6729
rect 544 6703 574 6729
rect 974 6703 1004 6729
rect 1060 6703 1090 6729
rect 458 6401 488 6503
rect 544 6401 574 6503
rect 458 6383 574 6401
rect 458 6349 499 6383
rect 533 6349 574 6383
rect 458 6331 574 6349
rect 974 6401 1004 6503
rect 1060 6401 1090 6503
rect 974 6383 1090 6401
rect 974 6349 1015 6383
rect 1049 6349 1090 6383
rect 974 6331 1090 6349
rect 458 5415 574 5433
rect 458 5381 499 5415
rect 533 5381 574 5415
rect 458 5363 574 5381
rect 458 5261 488 5363
rect 544 5261 574 5363
rect 974 5415 1090 5433
rect 974 5381 1015 5415
rect 1049 5381 1090 5415
rect 974 5363 1090 5381
rect 974 5261 1004 5363
rect 1060 5261 1090 5363
rect 458 5035 488 5061
rect 544 5035 574 5061
rect 974 5035 1004 5061
rect 1060 5035 1090 5061
rect 458 4255 574 4273
rect 458 4221 499 4255
rect 533 4221 574 4255
rect 458 4203 574 4221
rect 458 4101 488 4203
rect 544 4101 574 4203
rect 974 4255 1090 4273
rect 974 4221 1015 4255
rect 1049 4221 1090 4255
rect 974 4203 1090 4221
rect 974 4101 1004 4203
rect 1060 4101 1090 4203
rect 458 3675 488 3701
rect 544 3675 574 3701
rect 974 3675 1004 3701
rect 1060 3675 1090 3701
rect 458 3563 488 3589
rect 544 3563 574 3589
rect 974 3563 1004 3589
rect 1060 3563 1090 3589
rect 458 3125 488 3227
rect 544 3125 574 3227
rect 458 3107 574 3125
rect 458 3073 499 3107
rect 533 3073 574 3107
rect 458 3055 574 3073
rect 974 3125 1004 3227
rect 1060 3125 1090 3227
rect 974 3107 1090 3125
rect 974 3073 1015 3107
rect 1049 3073 1090 3107
rect 974 3055 1090 3073
rect 458 2491 574 2509
rect 458 2457 499 2491
rect 533 2457 574 2491
rect 458 2439 574 2457
rect 458 2337 488 2439
rect 544 2337 574 2439
rect 974 2491 1090 2509
rect 974 2457 1015 2491
rect 1049 2457 1090 2491
rect 974 2439 1090 2457
rect 974 2337 1004 2439
rect 1060 2337 1090 2439
rect 458 1975 488 2001
rect 544 1975 574 2001
rect 974 1975 1004 2001
rect 1060 1975 1090 2001
rect 458 1863 488 1889
rect 544 1863 574 1889
rect 974 1863 1004 1889
rect 1060 1863 1090 1889
rect 458 1425 488 1527
rect 544 1425 574 1527
rect 458 1407 574 1425
rect 458 1373 499 1407
rect 533 1373 574 1407
rect 458 1355 574 1373
rect 974 1425 1004 1527
rect 1060 1425 1090 1527
rect 974 1407 1090 1425
rect 974 1373 1015 1407
rect 1049 1373 1090 1407
rect 974 1355 1090 1373
<< polycont >>
rect 499 6349 533 6383
rect 1015 6349 1049 6383
rect 499 5381 533 5415
rect 1015 5381 1049 5415
rect 499 4221 533 4255
rect 1015 4221 1049 4255
rect 499 3073 533 3107
rect 1015 3073 1049 3107
rect 499 2457 533 2491
rect 1015 2457 1049 2491
rect 499 1373 533 1407
rect 1015 1373 1049 1407
<< locali >>
rect 413 7706 447 7714
rect 413 7634 447 7664
rect 413 7562 447 7596
rect 413 7494 447 7528
rect 413 7426 447 7456
rect 413 7376 447 7384
rect 499 7706 533 7714
rect 499 7634 533 7664
rect 499 7562 533 7596
rect 499 7494 533 7528
rect 499 7426 533 7456
rect 499 7376 533 7384
rect 585 7706 619 7714
rect 585 7634 619 7664
rect 585 7562 619 7596
rect 585 7494 619 7528
rect 585 7426 619 7456
rect 585 7376 619 7384
rect 671 7706 705 7714
rect 671 7634 705 7664
rect 671 7562 705 7596
rect 671 7494 705 7528
rect 671 7426 705 7456
rect 671 7376 705 7384
rect 757 7706 791 7714
rect 757 7634 791 7664
rect 757 7562 791 7596
rect 757 7494 791 7528
rect 757 7426 791 7456
rect 757 7376 791 7384
rect 843 7706 877 7714
rect 843 7634 877 7664
rect 843 7562 877 7596
rect 843 7494 877 7528
rect 843 7426 877 7456
rect 843 7376 877 7384
rect 929 7706 963 7714
rect 929 7634 963 7664
rect 929 7562 963 7596
rect 929 7494 963 7528
rect 929 7426 963 7456
rect 929 7376 963 7384
rect 1015 7706 1049 7714
rect 1015 7634 1049 7664
rect 1015 7562 1049 7596
rect 1015 7494 1049 7528
rect 1015 7426 1049 7456
rect 1015 7376 1049 7384
rect 1101 7706 1135 7714
rect 1101 7634 1135 7664
rect 1101 7562 1135 7596
rect 1101 7494 1135 7528
rect 1101 7426 1135 7456
rect 1101 7376 1135 7384
rect 413 6692 447 6704
rect 413 6620 447 6654
rect 413 6552 447 6586
rect 413 6502 447 6514
rect 499 6692 533 6704
rect 499 6620 533 6654
rect 499 6552 533 6586
rect 499 6502 533 6514
rect 585 6692 619 6704
rect 585 6620 619 6654
rect 585 6552 619 6586
rect 585 6502 619 6514
rect 929 6692 963 6704
rect 929 6620 963 6654
rect 929 6552 963 6586
rect 929 6502 963 6514
rect 1015 6692 1049 6704
rect 1015 6620 1049 6654
rect 1015 6552 1049 6586
rect 1015 6502 1049 6514
rect 1101 6692 1135 6704
rect 1101 6620 1135 6654
rect 1101 6552 1135 6586
rect 1101 6502 1135 6514
rect 482 6349 499 6383
rect 533 6349 550 6383
rect 998 6349 1015 6383
rect 1049 6349 1066 6383
rect 482 5381 499 5415
rect 533 5381 550 5415
rect 998 5381 1015 5415
rect 1049 5381 1066 5415
rect 413 5250 447 5262
rect 413 5178 447 5212
rect 413 5110 447 5144
rect 413 5060 447 5072
rect 499 5250 533 5262
rect 499 5178 533 5212
rect 499 5110 533 5144
rect 499 5060 533 5072
rect 585 5250 619 5262
rect 585 5178 619 5212
rect 585 5110 619 5144
rect 585 5060 619 5072
rect 929 5250 963 5262
rect 929 5178 963 5212
rect 929 5110 963 5144
rect 929 5060 963 5072
rect 1015 5250 1049 5262
rect 1015 5178 1049 5212
rect 1015 5110 1049 5144
rect 1015 5060 1049 5072
rect 1101 5250 1135 5262
rect 1101 5178 1135 5212
rect 1101 5110 1135 5144
rect 1101 5060 1135 5072
rect 482 4221 499 4255
rect 533 4221 550 4255
rect 998 4221 1015 4255
rect 1049 4221 1066 4255
rect 413 4088 447 4104
rect 413 4020 447 4028
rect 413 3952 447 3956
rect 413 3846 447 3850
rect 413 3774 447 3782
rect 413 3698 447 3714
rect 499 4088 533 4104
rect 499 4020 533 4028
rect 499 3952 533 3956
rect 499 3846 533 3850
rect 499 3774 533 3782
rect 499 3698 533 3714
rect 585 4088 619 4104
rect 585 4020 619 4028
rect 585 3952 619 3956
rect 585 3846 619 3850
rect 585 3774 619 3782
rect 585 3698 619 3714
rect 929 4088 963 4104
rect 929 4020 963 4028
rect 929 3952 963 3956
rect 929 3846 963 3850
rect 929 3774 963 3782
rect 929 3698 963 3714
rect 1015 4088 1049 4104
rect 1015 4020 1049 4028
rect 1015 3952 1049 3956
rect 1015 3846 1049 3850
rect 1015 3774 1049 3782
rect 1015 3698 1049 3714
rect 1101 4088 1135 4104
rect 1101 4020 1135 4028
rect 1101 3952 1135 3956
rect 1101 3846 1135 3850
rect 1101 3774 1135 3782
rect 1101 3698 1135 3714
rect 413 3556 447 3564
rect 413 3484 447 3514
rect 413 3412 447 3446
rect 413 3344 447 3378
rect 413 3276 447 3306
rect 413 3226 447 3234
rect 499 3556 533 3564
rect 499 3484 533 3514
rect 499 3412 533 3446
rect 499 3344 533 3378
rect 499 3276 533 3306
rect 499 3226 533 3234
rect 585 3556 619 3564
rect 585 3484 619 3514
rect 585 3412 619 3446
rect 585 3344 619 3378
rect 585 3276 619 3306
rect 585 3226 619 3234
rect 929 3556 963 3564
rect 929 3484 963 3514
rect 929 3412 963 3446
rect 929 3344 963 3378
rect 929 3276 963 3306
rect 929 3226 963 3234
rect 1015 3556 1049 3564
rect 1015 3484 1049 3514
rect 1015 3412 1049 3446
rect 1015 3344 1049 3378
rect 1015 3276 1049 3306
rect 1015 3226 1049 3234
rect 1101 3556 1135 3564
rect 1101 3484 1135 3514
rect 1101 3412 1135 3446
rect 1101 3344 1135 3378
rect 1101 3276 1135 3306
rect 1101 3226 1135 3234
rect 482 3073 499 3107
rect 533 3073 550 3107
rect 998 3073 1015 3107
rect 1049 3073 1066 3107
rect 482 2457 499 2491
rect 533 2457 550 2491
rect 998 2457 1015 2491
rect 1049 2457 1066 2491
rect 413 2330 447 2338
rect 413 2258 447 2288
rect 413 2186 447 2220
rect 413 2118 447 2152
rect 413 2050 447 2080
rect 413 2000 447 2008
rect 499 2330 533 2338
rect 499 2258 533 2288
rect 499 2186 533 2220
rect 499 2118 533 2152
rect 499 2050 533 2080
rect 499 2000 533 2008
rect 585 2330 619 2338
rect 585 2258 619 2288
rect 585 2186 619 2220
rect 585 2118 619 2152
rect 585 2050 619 2080
rect 585 2000 619 2008
rect 929 2330 963 2338
rect 929 2258 963 2288
rect 929 2186 963 2220
rect 929 2118 963 2152
rect 929 2050 963 2080
rect 929 2000 963 2008
rect 1015 2330 1049 2338
rect 1015 2258 1049 2288
rect 1015 2186 1049 2220
rect 1015 2118 1049 2152
rect 1015 2050 1049 2080
rect 1015 2000 1049 2008
rect 1101 2330 1135 2338
rect 1101 2258 1135 2288
rect 1101 2186 1135 2220
rect 1101 2118 1135 2152
rect 1101 2050 1135 2080
rect 1101 2000 1135 2008
rect 413 1856 447 1864
rect 413 1784 447 1814
rect 413 1712 447 1746
rect 413 1644 447 1678
rect 413 1576 447 1606
rect 413 1526 447 1534
rect 499 1856 533 1864
rect 499 1784 533 1814
rect 499 1712 533 1746
rect 499 1644 533 1678
rect 499 1576 533 1606
rect 499 1526 533 1534
rect 585 1856 619 1864
rect 585 1784 619 1814
rect 585 1712 619 1746
rect 585 1644 619 1678
rect 585 1576 619 1606
rect 585 1526 619 1534
rect 929 1856 963 1864
rect 929 1784 963 1814
rect 929 1712 963 1746
rect 929 1644 963 1678
rect 929 1576 963 1606
rect 929 1526 963 1534
rect 1015 1856 1049 1864
rect 1015 1784 1049 1814
rect 1015 1712 1049 1746
rect 1015 1644 1049 1678
rect 1015 1576 1049 1606
rect 1015 1526 1049 1534
rect 1101 1856 1135 1864
rect 1101 1784 1135 1814
rect 1101 1712 1135 1746
rect 1101 1644 1135 1678
rect 1101 1576 1135 1606
rect 1101 1526 1135 1534
rect 482 1373 499 1407
rect 533 1373 550 1407
rect 998 1373 1015 1407
rect 1049 1373 1066 1407
rect 413 582 447 598
rect 413 514 447 522
rect 413 446 447 450
rect 413 340 447 344
rect 413 268 447 276
rect 413 192 447 208
rect 499 582 533 598
rect 499 514 533 522
rect 499 446 533 450
rect 499 340 533 344
rect 499 268 533 276
rect 499 192 533 208
rect 585 582 619 598
rect 585 514 619 522
rect 585 446 619 450
rect 585 340 619 344
rect 585 268 619 276
rect 585 192 619 208
rect 671 582 705 598
rect 671 514 705 522
rect 671 446 705 450
rect 671 340 705 344
rect 671 268 705 276
rect 671 192 705 208
rect 757 582 791 598
rect 757 514 791 522
rect 757 446 791 450
rect 757 340 791 344
rect 757 268 791 276
rect 757 192 791 208
rect 843 582 877 598
rect 843 514 877 522
rect 843 446 877 450
rect 843 340 877 344
rect 843 268 877 276
rect 843 192 877 208
rect 929 582 963 598
rect 929 514 963 522
rect 929 446 963 450
rect 929 340 963 344
rect 929 268 963 276
rect 929 192 963 208
rect 1015 582 1049 598
rect 1015 514 1049 522
rect 1015 446 1049 450
rect 1015 340 1049 344
rect 1015 268 1049 276
rect 1015 192 1049 208
rect 1101 582 1135 598
rect 1101 514 1135 522
rect 1101 446 1135 450
rect 1101 340 1135 344
rect 1101 268 1135 276
rect 1101 192 1135 208
<< viali >>
rect 413 7698 447 7706
rect 413 7672 447 7698
rect 413 7630 447 7634
rect 413 7600 447 7630
rect 413 7528 447 7562
rect 413 7460 447 7490
rect 413 7456 447 7460
rect 413 7392 447 7418
rect 413 7384 447 7392
rect 499 7698 533 7706
rect 499 7672 533 7698
rect 499 7630 533 7634
rect 499 7600 533 7630
rect 499 7528 533 7562
rect 499 7460 533 7490
rect 499 7456 533 7460
rect 499 7392 533 7418
rect 499 7384 533 7392
rect 585 7698 619 7706
rect 585 7672 619 7698
rect 585 7630 619 7634
rect 585 7600 619 7630
rect 585 7528 619 7562
rect 585 7460 619 7490
rect 585 7456 619 7460
rect 585 7392 619 7418
rect 585 7384 619 7392
rect 671 7698 705 7706
rect 671 7672 705 7698
rect 671 7630 705 7634
rect 671 7600 705 7630
rect 671 7528 705 7562
rect 671 7460 705 7490
rect 671 7456 705 7460
rect 671 7392 705 7418
rect 671 7384 705 7392
rect 757 7698 791 7706
rect 757 7672 791 7698
rect 757 7630 791 7634
rect 757 7600 791 7630
rect 757 7528 791 7562
rect 757 7460 791 7490
rect 757 7456 791 7460
rect 757 7392 791 7418
rect 757 7384 791 7392
rect 843 7698 877 7706
rect 843 7672 877 7698
rect 843 7630 877 7634
rect 843 7600 877 7630
rect 843 7528 877 7562
rect 843 7460 877 7490
rect 843 7456 877 7460
rect 843 7392 877 7418
rect 843 7384 877 7392
rect 929 7698 963 7706
rect 929 7672 963 7698
rect 929 7630 963 7634
rect 929 7600 963 7630
rect 929 7528 963 7562
rect 929 7460 963 7490
rect 929 7456 963 7460
rect 929 7392 963 7418
rect 929 7384 963 7392
rect 1015 7698 1049 7706
rect 1015 7672 1049 7698
rect 1015 7630 1049 7634
rect 1015 7600 1049 7630
rect 1015 7528 1049 7562
rect 1015 7460 1049 7490
rect 1015 7456 1049 7460
rect 1015 7392 1049 7418
rect 1015 7384 1049 7392
rect 1101 7698 1135 7706
rect 1101 7672 1135 7698
rect 1101 7630 1135 7634
rect 1101 7600 1135 7630
rect 1101 7528 1135 7562
rect 1101 7460 1135 7490
rect 1101 7456 1135 7460
rect 1101 7392 1135 7418
rect 1101 7384 1135 7392
rect 413 6688 447 6692
rect 413 6658 447 6688
rect 413 6586 447 6620
rect 413 6518 447 6548
rect 413 6514 447 6518
rect 499 6688 533 6692
rect 499 6658 533 6688
rect 499 6586 533 6620
rect 499 6518 533 6548
rect 499 6514 533 6518
rect 585 6688 619 6692
rect 585 6658 619 6688
rect 585 6586 619 6620
rect 585 6518 619 6548
rect 585 6514 619 6518
rect 929 6688 963 6692
rect 929 6658 963 6688
rect 929 6586 963 6620
rect 929 6518 963 6548
rect 929 6514 963 6518
rect 1015 6688 1049 6692
rect 1015 6658 1049 6688
rect 1015 6586 1049 6620
rect 1015 6518 1049 6548
rect 1015 6514 1049 6518
rect 1101 6688 1135 6692
rect 1101 6658 1135 6688
rect 1101 6586 1135 6620
rect 1101 6518 1135 6548
rect 1101 6514 1135 6518
rect 499 6349 533 6383
rect 1015 6349 1049 6383
rect 499 5381 533 5415
rect 1015 5381 1049 5415
rect 413 5246 447 5250
rect 413 5216 447 5246
rect 413 5144 447 5178
rect 413 5076 447 5106
rect 413 5072 447 5076
rect 499 5246 533 5250
rect 499 5216 533 5246
rect 499 5144 533 5178
rect 499 5076 533 5106
rect 499 5072 533 5076
rect 585 5246 619 5250
rect 585 5216 619 5246
rect 585 5144 619 5178
rect 585 5076 619 5106
rect 585 5072 619 5076
rect 929 5246 963 5250
rect 929 5216 963 5246
rect 929 5144 963 5178
rect 929 5076 963 5106
rect 929 5072 963 5076
rect 1015 5246 1049 5250
rect 1015 5216 1049 5246
rect 1015 5144 1049 5178
rect 1015 5076 1049 5106
rect 1015 5072 1049 5076
rect 1101 5246 1135 5250
rect 1101 5216 1135 5246
rect 1101 5144 1135 5178
rect 1101 5076 1135 5106
rect 1101 5072 1135 5076
rect 499 4221 533 4255
rect 1015 4221 1049 4255
rect 413 4054 447 4062
rect 413 4028 447 4054
rect 413 3986 447 3990
rect 413 3956 447 3986
rect 413 3884 447 3918
rect 413 3816 447 3846
rect 413 3812 447 3816
rect 413 3748 447 3774
rect 413 3740 447 3748
rect 499 4054 533 4062
rect 499 4028 533 4054
rect 499 3986 533 3990
rect 499 3956 533 3986
rect 499 3884 533 3918
rect 499 3816 533 3846
rect 499 3812 533 3816
rect 499 3748 533 3774
rect 499 3740 533 3748
rect 585 4054 619 4062
rect 585 4028 619 4054
rect 585 3986 619 3990
rect 585 3956 619 3986
rect 585 3884 619 3918
rect 585 3816 619 3846
rect 585 3812 619 3816
rect 585 3748 619 3774
rect 585 3740 619 3748
rect 929 4054 963 4062
rect 929 4028 963 4054
rect 929 3986 963 3990
rect 929 3956 963 3986
rect 929 3884 963 3918
rect 929 3816 963 3846
rect 929 3812 963 3816
rect 929 3748 963 3774
rect 929 3740 963 3748
rect 1015 4054 1049 4062
rect 1015 4028 1049 4054
rect 1015 3986 1049 3990
rect 1015 3956 1049 3986
rect 1015 3884 1049 3918
rect 1015 3816 1049 3846
rect 1015 3812 1049 3816
rect 1015 3748 1049 3774
rect 1015 3740 1049 3748
rect 1101 4054 1135 4062
rect 1101 4028 1135 4054
rect 1101 3986 1135 3990
rect 1101 3956 1135 3986
rect 1101 3884 1135 3918
rect 1101 3816 1135 3846
rect 1101 3812 1135 3816
rect 1101 3748 1135 3774
rect 1101 3740 1135 3748
rect 413 3548 447 3556
rect 413 3522 447 3548
rect 413 3480 447 3484
rect 413 3450 447 3480
rect 413 3378 447 3412
rect 413 3310 447 3340
rect 413 3306 447 3310
rect 413 3242 447 3268
rect 413 3234 447 3242
rect 499 3548 533 3556
rect 499 3522 533 3548
rect 499 3480 533 3484
rect 499 3450 533 3480
rect 499 3378 533 3412
rect 499 3310 533 3340
rect 499 3306 533 3310
rect 499 3242 533 3268
rect 499 3234 533 3242
rect 585 3548 619 3556
rect 585 3522 619 3548
rect 585 3480 619 3484
rect 585 3450 619 3480
rect 585 3378 619 3412
rect 585 3310 619 3340
rect 585 3306 619 3310
rect 585 3242 619 3268
rect 585 3234 619 3242
rect 929 3548 963 3556
rect 929 3522 963 3548
rect 929 3480 963 3484
rect 929 3450 963 3480
rect 929 3378 963 3412
rect 929 3310 963 3340
rect 929 3306 963 3310
rect 929 3242 963 3268
rect 929 3234 963 3242
rect 1015 3548 1049 3556
rect 1015 3522 1049 3548
rect 1015 3480 1049 3484
rect 1015 3450 1049 3480
rect 1015 3378 1049 3412
rect 1015 3310 1049 3340
rect 1015 3306 1049 3310
rect 1015 3242 1049 3268
rect 1015 3234 1049 3242
rect 1101 3548 1135 3556
rect 1101 3522 1135 3548
rect 1101 3480 1135 3484
rect 1101 3450 1135 3480
rect 1101 3378 1135 3412
rect 1101 3310 1135 3340
rect 1101 3306 1135 3310
rect 1101 3242 1135 3268
rect 1101 3234 1135 3242
rect 499 3073 533 3107
rect 1015 3073 1049 3107
rect 499 2457 533 2491
rect 1015 2457 1049 2491
rect 413 2322 447 2330
rect 413 2296 447 2322
rect 413 2254 447 2258
rect 413 2224 447 2254
rect 413 2152 447 2186
rect 413 2084 447 2114
rect 413 2080 447 2084
rect 413 2016 447 2042
rect 413 2008 447 2016
rect 499 2322 533 2330
rect 499 2296 533 2322
rect 499 2254 533 2258
rect 499 2224 533 2254
rect 499 2152 533 2186
rect 499 2084 533 2114
rect 499 2080 533 2084
rect 499 2016 533 2042
rect 499 2008 533 2016
rect 585 2322 619 2330
rect 585 2296 619 2322
rect 585 2254 619 2258
rect 585 2224 619 2254
rect 585 2152 619 2186
rect 585 2084 619 2114
rect 585 2080 619 2084
rect 585 2016 619 2042
rect 585 2008 619 2016
rect 929 2322 963 2330
rect 929 2296 963 2322
rect 929 2254 963 2258
rect 929 2224 963 2254
rect 929 2152 963 2186
rect 929 2084 963 2114
rect 929 2080 963 2084
rect 929 2016 963 2042
rect 929 2008 963 2016
rect 1015 2322 1049 2330
rect 1015 2296 1049 2322
rect 1015 2254 1049 2258
rect 1015 2224 1049 2254
rect 1015 2152 1049 2186
rect 1015 2084 1049 2114
rect 1015 2080 1049 2084
rect 1015 2016 1049 2042
rect 1015 2008 1049 2016
rect 1101 2322 1135 2330
rect 1101 2296 1135 2322
rect 1101 2254 1135 2258
rect 1101 2224 1135 2254
rect 1101 2152 1135 2186
rect 1101 2084 1135 2114
rect 1101 2080 1135 2084
rect 1101 2016 1135 2042
rect 1101 2008 1135 2016
rect 413 1848 447 1856
rect 413 1822 447 1848
rect 413 1780 447 1784
rect 413 1750 447 1780
rect 413 1678 447 1712
rect 413 1610 447 1640
rect 413 1606 447 1610
rect 413 1542 447 1568
rect 413 1534 447 1542
rect 499 1848 533 1856
rect 499 1822 533 1848
rect 499 1780 533 1784
rect 499 1750 533 1780
rect 499 1678 533 1712
rect 499 1610 533 1640
rect 499 1606 533 1610
rect 499 1542 533 1568
rect 499 1534 533 1542
rect 585 1848 619 1856
rect 585 1822 619 1848
rect 585 1780 619 1784
rect 585 1750 619 1780
rect 585 1678 619 1712
rect 585 1610 619 1640
rect 585 1606 619 1610
rect 585 1542 619 1568
rect 585 1534 619 1542
rect 929 1848 963 1856
rect 929 1822 963 1848
rect 929 1780 963 1784
rect 929 1750 963 1780
rect 929 1678 963 1712
rect 929 1610 963 1640
rect 929 1606 963 1610
rect 929 1542 963 1568
rect 929 1534 963 1542
rect 1015 1848 1049 1856
rect 1015 1822 1049 1848
rect 1015 1780 1049 1784
rect 1015 1750 1049 1780
rect 1015 1678 1049 1712
rect 1015 1610 1049 1640
rect 1015 1606 1049 1610
rect 1015 1542 1049 1568
rect 1015 1534 1049 1542
rect 1101 1848 1135 1856
rect 1101 1822 1135 1848
rect 1101 1780 1135 1784
rect 1101 1750 1135 1780
rect 1101 1678 1135 1712
rect 1101 1610 1135 1640
rect 1101 1606 1135 1610
rect 1101 1542 1135 1568
rect 1101 1534 1135 1542
rect 499 1373 533 1407
rect 1015 1373 1049 1407
rect 413 548 447 556
rect 413 522 447 548
rect 413 480 447 484
rect 413 450 447 480
rect 413 378 447 412
rect 413 310 447 340
rect 413 306 447 310
rect 413 242 447 268
rect 413 234 447 242
rect 499 548 533 556
rect 499 522 533 548
rect 499 480 533 484
rect 499 450 533 480
rect 499 378 533 412
rect 499 310 533 340
rect 499 306 533 310
rect 499 242 533 268
rect 499 234 533 242
rect 585 548 619 556
rect 585 522 619 548
rect 585 480 619 484
rect 585 450 619 480
rect 585 378 619 412
rect 585 310 619 340
rect 585 306 619 310
rect 585 242 619 268
rect 585 234 619 242
rect 671 548 705 556
rect 671 522 705 548
rect 671 480 705 484
rect 671 450 705 480
rect 671 378 705 412
rect 671 310 705 340
rect 671 306 705 310
rect 671 242 705 268
rect 671 234 705 242
rect 757 548 791 556
rect 757 522 791 548
rect 757 480 791 484
rect 757 450 791 480
rect 757 378 791 412
rect 757 310 791 340
rect 757 306 791 310
rect 757 242 791 268
rect 757 234 791 242
rect 843 548 877 556
rect 843 522 877 548
rect 843 480 877 484
rect 843 450 877 480
rect 843 378 877 412
rect 843 310 877 340
rect 843 306 877 310
rect 843 242 877 268
rect 843 234 877 242
rect 929 548 963 556
rect 929 522 963 548
rect 929 480 963 484
rect 929 450 963 480
rect 929 378 963 412
rect 929 310 963 340
rect 929 306 963 310
rect 929 242 963 268
rect 929 234 963 242
rect 1015 548 1049 556
rect 1015 522 1049 548
rect 1015 480 1049 484
rect 1015 450 1049 480
rect 1015 378 1049 412
rect 1015 310 1049 340
rect 1015 306 1049 310
rect 1015 242 1049 268
rect 1015 234 1049 242
rect 1101 548 1135 556
rect 1101 522 1135 548
rect 1101 480 1135 484
rect 1101 450 1135 480
rect 1101 378 1135 412
rect 1101 310 1135 340
rect 1101 306 1135 310
rect 1101 242 1135 268
rect 1101 234 1135 242
<< metal1 >>
rect 404 7712 456 7718
rect 404 7634 456 7660
rect 404 7600 413 7634
rect 447 7600 456 7634
rect 404 7562 456 7600
rect 404 7528 413 7562
rect 447 7528 456 7562
rect 404 7490 456 7528
rect 404 7456 413 7490
rect 447 7456 456 7490
rect 404 7418 456 7456
rect 404 7384 413 7418
rect 447 7384 456 7418
rect 404 6692 456 7384
rect 490 7712 542 7718
rect 490 7634 542 7660
rect 490 7600 499 7634
rect 533 7600 542 7634
rect 490 7562 542 7600
rect 490 7528 499 7562
rect 533 7528 542 7562
rect 490 7490 542 7528
rect 490 7456 499 7490
rect 533 7456 542 7490
rect 490 7418 542 7456
rect 490 7384 499 7418
rect 533 7384 542 7418
rect 490 7372 542 7384
rect 576 7712 628 7718
rect 576 7634 628 7660
rect 576 7600 585 7634
rect 619 7600 628 7634
rect 576 7562 628 7600
rect 576 7528 585 7562
rect 619 7528 628 7562
rect 576 7490 628 7528
rect 576 7456 585 7490
rect 619 7456 628 7490
rect 576 7418 628 7456
rect 576 7384 585 7418
rect 619 7384 628 7418
rect 404 6658 413 6692
rect 447 6658 456 6692
rect 404 6620 456 6658
rect 404 6586 413 6620
rect 447 6586 456 6620
rect 404 6548 456 6586
rect 404 6514 413 6548
rect 447 6514 456 6548
rect 404 5250 456 6514
rect 490 6692 542 6704
rect 490 6658 499 6692
rect 533 6658 542 6692
rect 490 6620 542 6658
rect 490 6586 499 6620
rect 533 6586 542 6620
rect 490 6578 542 6586
rect 490 6514 499 6526
rect 533 6514 542 6526
rect 490 6502 542 6514
rect 576 6692 628 7384
rect 662 7712 714 7718
rect 662 7634 714 7660
rect 662 7600 671 7634
rect 705 7600 714 7634
rect 662 7562 714 7600
rect 662 7528 671 7562
rect 705 7528 714 7562
rect 662 7490 714 7528
rect 662 7456 671 7490
rect 705 7456 714 7490
rect 662 7418 714 7456
rect 662 7384 671 7418
rect 705 7384 714 7418
rect 662 7372 714 7384
rect 748 7712 800 7718
rect 748 7634 800 7660
rect 748 7600 757 7634
rect 791 7600 800 7634
rect 748 7562 800 7600
rect 748 7528 757 7562
rect 791 7528 800 7562
rect 748 7490 800 7528
rect 748 7456 757 7490
rect 791 7456 800 7490
rect 748 7418 800 7456
rect 748 7384 757 7418
rect 791 7384 800 7418
rect 748 7372 800 7384
rect 834 7712 886 7718
rect 834 7634 886 7660
rect 834 7600 843 7634
rect 877 7600 886 7634
rect 834 7562 886 7600
rect 834 7528 843 7562
rect 877 7528 886 7562
rect 834 7490 886 7528
rect 834 7456 843 7490
rect 877 7456 886 7490
rect 834 7418 886 7456
rect 834 7384 843 7418
rect 877 7384 886 7418
rect 834 7372 886 7384
rect 920 7712 972 7718
rect 920 7634 972 7660
rect 920 7600 929 7634
rect 963 7600 972 7634
rect 920 7562 972 7600
rect 920 7528 929 7562
rect 963 7528 972 7562
rect 920 7490 972 7528
rect 920 7456 929 7490
rect 963 7456 972 7490
rect 920 7418 972 7456
rect 920 7384 929 7418
rect 963 7384 972 7418
rect 576 6658 585 6692
rect 619 6658 628 6692
rect 576 6620 628 6658
rect 576 6586 585 6620
rect 619 6586 628 6620
rect 576 6548 628 6586
rect 576 6514 585 6548
rect 619 6514 628 6548
rect 490 6383 542 6395
rect 490 6349 499 6383
rect 533 6349 542 6383
rect 490 6200 542 6349
rect 490 6142 542 6148
rect 490 5444 542 5450
rect 490 5381 499 5392
rect 533 5381 542 5392
rect 490 5369 542 5381
rect 404 5216 413 5250
rect 447 5216 456 5250
rect 404 5178 456 5216
rect 404 5144 413 5178
rect 447 5144 456 5178
rect 404 5106 456 5144
rect 404 5072 413 5106
rect 447 5072 456 5106
rect 404 4062 456 5072
rect 490 5250 542 5262
rect 490 5216 499 5250
rect 533 5216 542 5250
rect 490 5178 542 5216
rect 490 5144 499 5178
rect 533 5144 542 5178
rect 490 5106 542 5144
rect 490 5072 499 5106
rect 533 5072 542 5106
rect 490 5066 542 5072
rect 490 5008 542 5014
rect 576 5250 628 6514
rect 576 5216 585 5250
rect 619 5216 628 5250
rect 576 5178 628 5216
rect 576 5144 585 5178
rect 619 5144 628 5178
rect 576 5106 628 5144
rect 576 5072 585 5106
rect 619 5072 628 5106
rect 490 4310 542 4316
rect 490 4255 542 4258
rect 490 4221 499 4255
rect 533 4221 542 4255
rect 490 4209 542 4221
rect 404 4028 413 4062
rect 447 4028 456 4062
rect 404 3990 456 4028
rect 404 3956 413 3990
rect 447 3956 456 3990
rect 404 3918 456 3956
rect 404 3884 413 3918
rect 447 3884 456 3918
rect 404 3846 456 3884
rect 404 3812 413 3846
rect 447 3812 456 3846
rect 404 3774 456 3812
rect 404 3740 413 3774
rect 447 3740 456 3774
rect 404 3728 456 3740
rect 490 4062 542 4074
rect 490 4028 499 4062
rect 533 4028 542 4062
rect 490 3990 542 4028
rect 490 3956 499 3990
rect 533 3956 542 3990
rect 490 3918 542 3956
rect 490 3884 499 3918
rect 533 3884 542 3918
rect 490 3846 542 3884
rect 490 3812 499 3846
rect 533 3812 542 3846
rect 490 3774 542 3812
rect 490 3740 499 3774
rect 533 3740 542 3774
rect 404 3556 456 3568
rect 404 3522 413 3556
rect 447 3522 456 3556
rect 404 3484 456 3522
rect 404 3450 413 3484
rect 447 3450 456 3484
rect 404 3412 456 3450
rect 404 3378 413 3412
rect 447 3378 456 3412
rect 404 3340 456 3378
rect 404 3306 413 3340
rect 447 3306 456 3340
rect 404 3302 456 3306
rect 404 3234 413 3250
rect 447 3234 456 3250
rect 404 2330 456 3234
rect 490 3556 542 3740
rect 576 4062 628 5072
rect 576 4028 585 4062
rect 619 4028 628 4062
rect 576 3990 628 4028
rect 576 3956 585 3990
rect 619 3956 628 3990
rect 576 3918 628 3956
rect 576 3884 585 3918
rect 619 3884 628 3918
rect 576 3846 628 3884
rect 576 3812 585 3846
rect 619 3812 628 3846
rect 576 3774 628 3812
rect 576 3740 585 3774
rect 619 3740 628 3774
rect 576 3728 628 3740
rect 920 6692 972 7384
rect 1006 7712 1058 7718
rect 1006 7634 1058 7660
rect 1006 7600 1015 7634
rect 1049 7600 1058 7634
rect 1006 7562 1058 7600
rect 1006 7528 1015 7562
rect 1049 7528 1058 7562
rect 1006 7490 1058 7528
rect 1006 7456 1015 7490
rect 1049 7456 1058 7490
rect 1006 7418 1058 7456
rect 1006 7384 1015 7418
rect 1049 7384 1058 7418
rect 1006 7372 1058 7384
rect 1092 7712 1144 7718
rect 1092 7634 1144 7660
rect 1092 7600 1101 7634
rect 1135 7600 1144 7634
rect 1092 7562 1144 7600
rect 1092 7528 1101 7562
rect 1135 7528 1144 7562
rect 1092 7490 1144 7528
rect 1092 7456 1101 7490
rect 1135 7456 1144 7490
rect 1092 7418 1144 7456
rect 1092 7384 1101 7418
rect 1135 7384 1144 7418
rect 920 6658 929 6692
rect 963 6658 972 6692
rect 920 6620 972 6658
rect 920 6586 929 6620
rect 963 6586 972 6620
rect 920 6548 972 6586
rect 920 6514 929 6548
rect 963 6514 972 6548
rect 920 5250 972 6514
rect 1006 6692 1058 6704
rect 1006 6658 1015 6692
rect 1049 6658 1058 6692
rect 1006 6620 1058 6658
rect 1006 6586 1015 6620
rect 1049 6586 1058 6620
rect 1006 6578 1058 6586
rect 1006 6514 1015 6526
rect 1049 6514 1058 6526
rect 1006 6502 1058 6514
rect 1092 6692 1144 7384
rect 1092 6658 1101 6692
rect 1135 6658 1144 6692
rect 1092 6620 1144 6658
rect 1092 6586 1101 6620
rect 1135 6586 1144 6620
rect 1092 6548 1144 6586
rect 1092 6514 1101 6548
rect 1135 6514 1144 6548
rect 1006 6383 1058 6395
rect 1006 6349 1015 6383
rect 1049 6349 1058 6383
rect 1006 6200 1058 6349
rect 1006 6142 1058 6148
rect 1006 5444 1058 5450
rect 1006 5381 1015 5392
rect 1049 5381 1058 5392
rect 1006 5369 1058 5381
rect 920 5216 929 5250
rect 963 5216 972 5250
rect 920 5178 972 5216
rect 920 5144 929 5178
rect 963 5144 972 5178
rect 920 5106 972 5144
rect 920 5072 929 5106
rect 963 5072 972 5106
rect 920 4062 972 5072
rect 1006 5250 1058 5262
rect 1006 5216 1015 5250
rect 1049 5216 1058 5250
rect 1006 5178 1058 5216
rect 1006 5144 1015 5178
rect 1049 5144 1058 5178
rect 1006 5106 1058 5144
rect 1006 5072 1015 5106
rect 1049 5072 1058 5106
rect 1006 5066 1058 5072
rect 1006 5008 1058 5014
rect 1092 5250 1144 6514
rect 1092 5216 1101 5250
rect 1135 5216 1144 5250
rect 1092 5178 1144 5216
rect 1092 5144 1101 5178
rect 1135 5144 1144 5178
rect 1092 5106 1144 5144
rect 1092 5072 1101 5106
rect 1135 5072 1144 5106
rect 1006 4310 1058 4316
rect 1006 4255 1058 4258
rect 1006 4221 1015 4255
rect 1049 4221 1058 4255
rect 1006 4209 1058 4221
rect 920 4028 929 4062
rect 963 4028 972 4062
rect 920 3990 972 4028
rect 920 3956 929 3990
rect 963 3956 972 3990
rect 920 3918 972 3956
rect 920 3884 929 3918
rect 963 3884 972 3918
rect 920 3846 972 3884
rect 920 3812 929 3846
rect 963 3812 972 3846
rect 920 3774 972 3812
rect 920 3740 929 3774
rect 963 3740 972 3774
rect 920 3728 972 3740
rect 1006 4062 1058 4074
rect 1006 4028 1015 4062
rect 1049 4028 1058 4062
rect 1006 3990 1058 4028
rect 1006 3956 1015 3990
rect 1049 3956 1058 3990
rect 1006 3918 1058 3956
rect 1006 3884 1015 3918
rect 1049 3884 1058 3918
rect 1006 3869 1058 3884
rect 1006 3812 1015 3817
rect 1049 3812 1058 3817
rect 1006 3774 1058 3812
rect 1006 3740 1015 3774
rect 1049 3740 1058 3774
rect 490 3522 499 3556
rect 533 3522 542 3556
rect 490 3491 542 3522
rect 490 3412 542 3439
rect 490 3378 499 3412
rect 533 3378 542 3412
rect 490 3340 542 3378
rect 490 3306 499 3340
rect 533 3306 542 3340
rect 490 3268 542 3306
rect 490 3234 499 3268
rect 533 3234 542 3268
rect 490 3222 542 3234
rect 576 3556 628 3568
rect 576 3522 585 3556
rect 619 3522 628 3556
rect 576 3484 628 3522
rect 576 3450 585 3484
rect 619 3450 628 3484
rect 576 3412 628 3450
rect 576 3378 585 3412
rect 619 3378 628 3412
rect 576 3340 628 3378
rect 576 3306 585 3340
rect 619 3306 628 3340
rect 576 3302 628 3306
rect 576 3234 585 3250
rect 619 3234 628 3250
rect 490 3113 542 3119
rect 490 3055 542 3061
rect 490 2735 542 2741
rect 490 2491 542 2683
rect 490 2457 499 2491
rect 533 2457 542 2491
rect 490 2445 542 2457
rect 404 2296 413 2330
rect 447 2296 456 2330
rect 404 2258 456 2296
rect 404 2224 413 2258
rect 447 2224 456 2258
rect 404 2186 456 2224
rect 404 2152 413 2186
rect 447 2152 456 2186
rect 404 2114 456 2152
rect 404 2080 413 2114
rect 447 2080 456 2114
rect 404 2042 456 2080
rect 404 2008 413 2042
rect 447 2008 456 2042
rect 404 1996 456 2008
rect 490 2330 542 2342
rect 490 2296 499 2330
rect 533 2296 542 2330
rect 490 2258 542 2296
rect 490 2224 499 2258
rect 533 2224 542 2258
rect 490 2186 542 2224
rect 490 2152 499 2186
rect 533 2152 542 2186
rect 490 2114 542 2152
rect 490 2105 499 2114
rect 533 2105 542 2114
rect 490 2042 542 2053
rect 490 2008 499 2042
rect 533 2008 542 2042
rect 404 1856 456 1868
rect 404 1822 413 1856
rect 447 1822 456 1856
rect 404 1784 456 1822
rect 404 1750 413 1784
rect 447 1750 456 1784
rect 404 1712 456 1750
rect 404 1678 413 1712
rect 447 1678 456 1712
rect 404 1640 456 1678
rect 404 1606 413 1640
rect 447 1606 456 1640
rect 404 1568 456 1606
rect 404 1534 413 1568
rect 447 1534 456 1568
rect 404 556 456 1534
rect 490 1856 542 2008
rect 576 2330 628 3234
rect 576 2296 585 2330
rect 619 2296 628 2330
rect 576 2258 628 2296
rect 576 2224 585 2258
rect 619 2224 628 2258
rect 576 2186 628 2224
rect 576 2152 585 2186
rect 619 2152 628 2186
rect 576 2114 628 2152
rect 576 2080 585 2114
rect 619 2080 628 2114
rect 576 2042 628 2080
rect 576 2008 585 2042
rect 619 2008 628 2042
rect 576 1996 628 2008
rect 920 3556 972 3568
rect 920 3522 929 3556
rect 963 3522 972 3556
rect 920 3484 972 3522
rect 920 3450 929 3484
rect 963 3450 972 3484
rect 920 3412 972 3450
rect 920 3378 929 3412
rect 963 3378 972 3412
rect 920 3340 972 3378
rect 920 3306 929 3340
rect 963 3306 972 3340
rect 920 3302 972 3306
rect 920 3234 929 3250
rect 963 3234 972 3250
rect 920 2330 972 3234
rect 1006 3556 1058 3740
rect 1092 4062 1144 5072
rect 1092 4028 1101 4062
rect 1135 4028 1144 4062
rect 1092 3990 1144 4028
rect 1092 3956 1101 3990
rect 1135 3956 1144 3990
rect 1092 3918 1144 3956
rect 1092 3884 1101 3918
rect 1135 3884 1144 3918
rect 1092 3846 1144 3884
rect 1092 3812 1101 3846
rect 1135 3812 1144 3846
rect 1092 3774 1144 3812
rect 1092 3740 1101 3774
rect 1135 3740 1144 3774
rect 1092 3728 1144 3740
rect 1006 3522 1015 3556
rect 1049 3522 1058 3556
rect 1006 3484 1058 3522
rect 1006 3450 1015 3484
rect 1049 3450 1058 3484
rect 1006 3412 1058 3450
rect 1006 3378 1015 3412
rect 1049 3378 1058 3412
rect 1006 3340 1058 3378
rect 1006 3306 1015 3340
rect 1049 3306 1058 3340
rect 1006 3268 1058 3306
rect 1006 3234 1015 3268
rect 1049 3234 1058 3268
rect 1006 3222 1058 3234
rect 1092 3556 1144 3568
rect 1092 3522 1101 3556
rect 1135 3522 1144 3556
rect 1092 3484 1144 3522
rect 1092 3450 1101 3484
rect 1135 3450 1144 3484
rect 1092 3412 1144 3450
rect 1092 3378 1101 3412
rect 1135 3378 1144 3412
rect 1092 3340 1144 3378
rect 1092 3306 1101 3340
rect 1135 3306 1144 3340
rect 1092 3302 1144 3306
rect 1092 3234 1101 3250
rect 1135 3234 1144 3250
rect 1006 3113 1058 3119
rect 1006 3055 1058 3061
rect 1006 2546 1058 2741
rect 1006 2491 1058 2494
rect 1006 2457 1015 2491
rect 1049 2457 1058 2491
rect 1006 2445 1058 2457
rect 920 2296 929 2330
rect 963 2296 972 2330
rect 920 2258 972 2296
rect 920 2224 929 2258
rect 963 2224 972 2258
rect 920 2186 972 2224
rect 920 2152 929 2186
rect 963 2152 972 2186
rect 920 2114 972 2152
rect 920 2080 929 2114
rect 963 2080 972 2114
rect 920 2042 972 2080
rect 920 2008 929 2042
rect 963 2008 972 2042
rect 920 1996 972 2008
rect 1006 2330 1058 2342
rect 1006 2296 1015 2330
rect 1049 2296 1058 2330
rect 1006 2258 1058 2296
rect 1006 2224 1015 2258
rect 1049 2224 1058 2258
rect 1006 2186 1058 2224
rect 1006 2152 1015 2186
rect 1049 2152 1058 2186
rect 1006 2114 1058 2152
rect 1006 2105 1015 2114
rect 1049 2105 1058 2114
rect 1006 2042 1058 2053
rect 1006 2008 1015 2042
rect 1049 2008 1058 2042
rect 490 1822 499 1856
rect 533 1822 542 1856
rect 490 1784 542 1822
rect 490 1750 499 1784
rect 533 1750 542 1784
rect 490 1712 542 1750
rect 490 1678 499 1712
rect 533 1678 542 1712
rect 490 1640 542 1678
rect 490 1606 499 1640
rect 533 1606 542 1640
rect 490 1568 542 1606
rect 490 1534 499 1568
rect 533 1534 542 1568
rect 490 1522 542 1534
rect 576 1856 628 1868
rect 576 1822 585 1856
rect 619 1822 628 1856
rect 576 1784 628 1822
rect 576 1750 585 1784
rect 619 1750 628 1784
rect 576 1712 628 1750
rect 576 1678 585 1712
rect 619 1678 628 1712
rect 576 1640 628 1678
rect 576 1606 585 1640
rect 619 1606 628 1640
rect 576 1568 628 1606
rect 576 1534 585 1568
rect 619 1534 628 1568
rect 490 1412 542 1419
rect 490 1354 542 1360
rect 404 530 413 556
rect 447 530 456 556
rect 404 450 413 478
rect 447 450 456 478
rect 404 412 456 450
rect 404 378 413 412
rect 447 378 456 412
rect 404 340 456 378
rect 404 306 413 340
rect 447 306 456 340
rect 404 268 456 306
rect 404 234 413 268
rect 447 234 456 268
rect 404 222 456 234
rect 490 556 542 568
rect 490 530 499 556
rect 533 530 542 556
rect 490 450 499 478
rect 533 450 542 478
rect 490 412 542 450
rect 490 378 499 412
rect 533 378 542 412
rect 490 340 542 378
rect 490 306 499 340
rect 533 306 542 340
rect 490 268 542 306
rect 490 234 499 268
rect 533 234 542 268
rect 490 222 542 234
rect 576 556 628 1534
rect 920 1856 972 1868
rect 920 1822 929 1856
rect 963 1822 972 1856
rect 920 1784 972 1822
rect 920 1750 929 1784
rect 963 1750 972 1784
rect 920 1712 972 1750
rect 920 1678 929 1712
rect 963 1678 972 1712
rect 920 1640 972 1678
rect 920 1606 929 1640
rect 963 1606 972 1640
rect 920 1568 972 1606
rect 920 1534 929 1568
rect 963 1534 972 1568
rect 576 530 585 556
rect 619 530 628 556
rect 576 450 585 478
rect 619 450 628 478
rect 576 412 628 450
rect 576 378 585 412
rect 619 378 628 412
rect 576 340 628 378
rect 576 306 585 340
rect 619 306 628 340
rect 576 268 628 306
rect 576 234 585 268
rect 619 234 628 268
rect 576 222 628 234
rect 662 556 714 568
rect 662 530 671 556
rect 705 530 714 556
rect 662 450 671 478
rect 705 450 714 478
rect 662 412 714 450
rect 662 378 671 412
rect 705 378 714 412
rect 662 340 714 378
rect 662 306 671 340
rect 705 306 714 340
rect 662 268 714 306
rect 662 234 671 268
rect 705 234 714 268
rect 662 222 714 234
rect 748 556 800 568
rect 748 530 757 556
rect 791 530 800 556
rect 748 450 757 478
rect 791 450 800 478
rect 748 412 800 450
rect 748 378 757 412
rect 791 378 800 412
rect 748 340 800 378
rect 748 306 757 340
rect 791 306 800 340
rect 748 268 800 306
rect 748 234 757 268
rect 791 234 800 268
rect 748 222 800 234
rect 834 556 886 568
rect 834 530 843 556
rect 877 530 886 556
rect 834 450 843 478
rect 877 450 886 478
rect 834 412 886 450
rect 834 378 843 412
rect 877 378 886 412
rect 834 340 886 378
rect 834 306 843 340
rect 877 306 886 340
rect 834 268 886 306
rect 834 234 843 268
rect 877 234 886 268
rect 834 222 886 234
rect 920 556 972 1534
rect 1006 1856 1058 2008
rect 1092 2330 1144 3234
rect 1092 2296 1101 2330
rect 1135 2296 1144 2330
rect 1092 2258 1144 2296
rect 1092 2224 1101 2258
rect 1135 2224 1144 2258
rect 1092 2186 1144 2224
rect 1092 2152 1101 2186
rect 1135 2152 1144 2186
rect 1092 2114 1144 2152
rect 1092 2080 1101 2114
rect 1135 2080 1144 2114
rect 1092 2042 1144 2080
rect 1092 2008 1101 2042
rect 1135 2008 1144 2042
rect 1092 1996 1144 2008
rect 1006 1822 1015 1856
rect 1049 1822 1058 1856
rect 1006 1784 1058 1822
rect 1006 1750 1015 1784
rect 1049 1750 1058 1784
rect 1006 1712 1058 1750
rect 1006 1678 1015 1712
rect 1049 1678 1058 1712
rect 1006 1640 1058 1678
rect 1006 1606 1015 1640
rect 1049 1606 1058 1640
rect 1006 1568 1058 1606
rect 1006 1534 1015 1568
rect 1049 1534 1058 1568
rect 1006 1522 1058 1534
rect 1092 1856 1144 1868
rect 1092 1822 1101 1856
rect 1135 1822 1144 1856
rect 1092 1784 1144 1822
rect 1092 1750 1101 1784
rect 1135 1750 1144 1784
rect 1092 1712 1144 1750
rect 1092 1678 1101 1712
rect 1135 1678 1144 1712
rect 1092 1640 1144 1678
rect 1092 1606 1101 1640
rect 1135 1606 1144 1640
rect 1092 1568 1144 1606
rect 1092 1534 1101 1568
rect 1135 1534 1144 1568
rect 1006 1412 1058 1419
rect 1006 1354 1058 1360
rect 920 530 929 556
rect 963 530 972 556
rect 920 450 929 478
rect 963 450 972 478
rect 920 412 972 450
rect 920 378 929 412
rect 963 378 972 412
rect 920 340 972 378
rect 920 306 929 340
rect 963 306 972 340
rect 920 268 972 306
rect 920 234 929 268
rect 963 234 972 268
rect 920 222 972 234
rect 1006 556 1058 568
rect 1006 530 1015 556
rect 1049 530 1058 556
rect 1006 450 1015 478
rect 1049 450 1058 478
rect 1006 412 1058 450
rect 1006 378 1015 412
rect 1049 378 1058 412
rect 1006 340 1058 378
rect 1006 306 1015 340
rect 1049 306 1058 340
rect 1006 268 1058 306
rect 1006 234 1015 268
rect 1049 234 1058 268
rect 1006 222 1058 234
rect 1092 556 1144 1534
rect 1092 530 1101 556
rect 1135 530 1144 556
rect 1092 450 1101 478
rect 1135 450 1144 478
rect 1092 412 1144 450
rect 1092 378 1101 412
rect 1135 378 1144 412
rect 1092 340 1144 378
rect 1092 306 1101 340
rect 1135 306 1144 340
rect 1092 268 1144 306
rect 1092 234 1101 268
rect 1135 234 1144 268
rect 1092 222 1144 234
<< via1 >>
rect 404 7706 456 7712
rect 404 7672 413 7706
rect 413 7672 447 7706
rect 447 7672 456 7706
rect 404 7660 456 7672
rect 490 7706 542 7712
rect 490 7672 499 7706
rect 499 7672 533 7706
rect 533 7672 542 7706
rect 490 7660 542 7672
rect 576 7706 628 7712
rect 576 7672 585 7706
rect 585 7672 619 7706
rect 619 7672 628 7706
rect 576 7660 628 7672
rect 490 6548 542 6578
rect 490 6526 499 6548
rect 499 6526 533 6548
rect 533 6526 542 6548
rect 662 7706 714 7712
rect 662 7672 671 7706
rect 671 7672 705 7706
rect 705 7672 714 7706
rect 662 7660 714 7672
rect 748 7706 800 7712
rect 748 7672 757 7706
rect 757 7672 791 7706
rect 791 7672 800 7706
rect 748 7660 800 7672
rect 834 7706 886 7712
rect 834 7672 843 7706
rect 843 7672 877 7706
rect 877 7672 886 7706
rect 834 7660 886 7672
rect 920 7706 972 7712
rect 920 7672 929 7706
rect 929 7672 963 7706
rect 963 7672 972 7706
rect 920 7660 972 7672
rect 490 6148 542 6200
rect 490 5415 542 5444
rect 490 5392 499 5415
rect 499 5392 533 5415
rect 533 5392 542 5415
rect 490 5014 542 5066
rect 490 4258 542 4310
rect 404 3268 456 3302
rect 404 3250 413 3268
rect 413 3250 447 3268
rect 447 3250 456 3268
rect 1006 7706 1058 7712
rect 1006 7672 1015 7706
rect 1015 7672 1049 7706
rect 1049 7672 1058 7706
rect 1006 7660 1058 7672
rect 1092 7706 1144 7712
rect 1092 7672 1101 7706
rect 1101 7672 1135 7706
rect 1135 7672 1144 7706
rect 1092 7660 1144 7672
rect 1006 6548 1058 6578
rect 1006 6526 1015 6548
rect 1015 6526 1049 6548
rect 1049 6526 1058 6548
rect 1006 6148 1058 6200
rect 1006 5415 1058 5444
rect 1006 5392 1015 5415
rect 1015 5392 1049 5415
rect 1049 5392 1058 5415
rect 1006 5014 1058 5066
rect 1006 4258 1058 4310
rect 1006 3846 1058 3869
rect 1006 3817 1015 3846
rect 1015 3817 1049 3846
rect 1049 3817 1058 3846
rect 490 3484 542 3491
rect 490 3450 499 3484
rect 499 3450 533 3484
rect 533 3450 542 3484
rect 490 3439 542 3450
rect 576 3268 628 3302
rect 576 3250 585 3268
rect 585 3250 619 3268
rect 619 3250 628 3268
rect 490 3107 542 3113
rect 490 3073 499 3107
rect 499 3073 533 3107
rect 533 3073 542 3107
rect 490 3061 542 3073
rect 490 2683 542 2735
rect 490 2080 499 2105
rect 499 2080 533 2105
rect 533 2080 542 2105
rect 490 2053 542 2080
rect 920 3268 972 3302
rect 920 3250 929 3268
rect 929 3250 963 3268
rect 963 3250 972 3268
rect 1092 3268 1144 3302
rect 1092 3250 1101 3268
rect 1101 3250 1135 3268
rect 1135 3250 1144 3268
rect 1006 3107 1058 3113
rect 1006 3073 1015 3107
rect 1015 3073 1049 3107
rect 1049 3073 1058 3107
rect 1006 3061 1058 3073
rect 1006 2494 1058 2546
rect 1006 2080 1015 2105
rect 1015 2080 1049 2105
rect 1049 2080 1058 2105
rect 1006 2053 1058 2080
rect 490 1407 542 1412
rect 490 1373 499 1407
rect 499 1373 533 1407
rect 533 1373 542 1407
rect 490 1360 542 1373
rect 404 522 413 530
rect 413 522 447 530
rect 447 522 456 530
rect 404 484 456 522
rect 404 478 413 484
rect 413 478 447 484
rect 447 478 456 484
rect 490 522 499 530
rect 499 522 533 530
rect 533 522 542 530
rect 490 484 542 522
rect 490 478 499 484
rect 499 478 533 484
rect 533 478 542 484
rect 576 522 585 530
rect 585 522 619 530
rect 619 522 628 530
rect 576 484 628 522
rect 576 478 585 484
rect 585 478 619 484
rect 619 478 628 484
rect 662 522 671 530
rect 671 522 705 530
rect 705 522 714 530
rect 662 484 714 522
rect 662 478 671 484
rect 671 478 705 484
rect 705 478 714 484
rect 748 522 757 530
rect 757 522 791 530
rect 791 522 800 530
rect 748 484 800 522
rect 748 478 757 484
rect 757 478 791 484
rect 791 478 800 484
rect 834 522 843 530
rect 843 522 877 530
rect 877 522 886 530
rect 834 484 886 522
rect 834 478 843 484
rect 843 478 877 484
rect 877 478 886 484
rect 1006 1407 1058 1412
rect 1006 1373 1015 1407
rect 1015 1373 1049 1407
rect 1049 1373 1058 1407
rect 1006 1360 1058 1373
rect 920 522 929 530
rect 929 522 963 530
rect 963 522 972 530
rect 920 484 972 522
rect 920 478 929 484
rect 929 478 963 484
rect 963 478 972 484
rect 1006 522 1015 530
rect 1015 522 1049 530
rect 1049 522 1058 530
rect 1006 484 1058 522
rect 1006 478 1015 484
rect 1015 478 1049 484
rect 1049 478 1058 484
rect 1092 522 1101 530
rect 1101 522 1135 530
rect 1135 522 1144 530
rect 1092 484 1144 522
rect 1092 478 1101 484
rect 1101 478 1135 484
rect 1135 478 1144 484
<< metal2 >>
rect 398 7712 1150 7714
rect 398 7660 404 7712
rect 456 7660 490 7712
rect 542 7660 576 7712
rect 628 7660 662 7712
rect 714 7660 748 7712
rect 800 7660 834 7712
rect 886 7660 920 7712
rect 972 7660 1006 7712
rect 1058 7660 1092 7712
rect 1144 7660 1150 7712
rect 398 7658 1150 7660
rect 484 6578 660 6580
rect 484 6526 490 6578
rect 542 6526 660 6578
rect 484 6524 660 6526
rect 716 6524 725 6580
rect 823 6524 832 6580
rect 888 6578 1064 6580
rect 888 6526 1006 6578
rect 1058 6526 1064 6578
rect 888 6524 1064 6526
rect 350 6146 359 6202
rect 415 6200 548 6202
rect 415 6148 490 6200
rect 542 6148 548 6200
rect 415 6146 548 6148
rect 1000 6200 1133 6202
rect 1000 6148 1006 6200
rect 1058 6148 1133 6200
rect 1000 6146 1133 6148
rect 1189 6146 1198 6202
rect 350 5390 359 5446
rect 415 5444 548 5446
rect 415 5392 490 5444
rect 542 5392 548 5444
rect 415 5390 548 5392
rect 1000 5444 1133 5446
rect 1000 5392 1006 5444
rect 1058 5392 1133 5444
rect 1000 5390 1133 5392
rect 1189 5390 1198 5446
rect 479 5012 488 5068
rect 544 5012 553 5068
rect 995 5012 1004 5068
rect 1060 5012 1069 5068
rect 479 4256 488 4312
rect 544 4256 553 4312
rect 995 4256 1004 4312
rect 1060 4256 1069 4312
rect 479 3815 488 3871
rect 544 3869 1064 3871
rect 544 3817 1006 3869
rect 1058 3817 1064 3869
rect 544 3815 1064 3817
rect 484 3491 1004 3493
rect 484 3439 490 3491
rect 542 3439 1004 3491
rect 484 3437 1004 3439
rect 1060 3437 1069 3493
rect 398 3302 660 3304
rect 398 3250 404 3302
rect 456 3250 576 3302
rect 628 3250 660 3302
rect 398 3248 660 3250
rect 716 3248 725 3304
rect 823 3248 832 3304
rect 888 3302 1150 3304
rect 888 3250 920 3302
rect 972 3250 1092 3302
rect 1144 3250 1150 3302
rect 888 3248 1150 3250
rect 479 3059 488 3115
rect 544 3059 553 3115
rect 995 3059 1004 3115
rect 1060 3059 1069 3115
rect 484 2735 1064 2737
rect 484 2683 490 2735
rect 542 2683 1064 2735
rect 484 2681 1064 2683
rect 484 2546 1064 2548
rect 484 2494 1006 2546
rect 1058 2494 1064 2546
rect 484 2492 1064 2494
rect 484 2105 1064 2107
rect 484 2053 490 2105
rect 542 2053 1006 2105
rect 1058 2053 1064 2105
rect 484 2051 1064 2053
rect 350 1358 359 1414
rect 415 1412 1133 1414
rect 415 1360 490 1412
rect 542 1360 1006 1412
rect 1058 1360 1133 1412
rect 415 1358 1133 1360
rect 1189 1358 1198 1414
rect 398 530 1150 532
rect 398 478 404 530
rect 456 478 490 530
rect 542 478 576 530
rect 628 478 662 530
rect 714 478 748 530
rect 800 478 834 530
rect 886 478 920 530
rect 972 478 1006 530
rect 1058 478 1092 530
rect 1144 478 1150 530
rect 398 476 1150 478
<< via2 >>
rect 660 6524 716 6580
rect 832 6524 888 6580
rect 359 6146 415 6202
rect 1133 6146 1189 6202
rect 359 5390 415 5446
rect 1133 5390 1189 5446
rect 488 5066 544 5068
rect 488 5014 490 5066
rect 490 5014 542 5066
rect 542 5014 544 5066
rect 488 5012 544 5014
rect 1004 5066 1060 5068
rect 1004 5014 1006 5066
rect 1006 5014 1058 5066
rect 1058 5014 1060 5066
rect 1004 5012 1060 5014
rect 488 4310 544 4312
rect 488 4258 490 4310
rect 490 4258 542 4310
rect 542 4258 544 4310
rect 488 4256 544 4258
rect 1004 4310 1060 4312
rect 1004 4258 1006 4310
rect 1006 4258 1058 4310
rect 1058 4258 1060 4310
rect 1004 4256 1060 4258
rect 488 3815 544 3871
rect 1004 3437 1060 3493
rect 660 3248 716 3304
rect 832 3248 888 3304
rect 488 3113 544 3115
rect 488 3061 490 3113
rect 490 3061 542 3113
rect 542 3061 544 3113
rect 488 3059 544 3061
rect 1004 3113 1060 3115
rect 1004 3061 1006 3113
rect 1006 3061 1058 3113
rect 1058 3061 1060 3113
rect 1004 3059 1060 3061
rect 359 1358 415 1414
rect 1133 1358 1189 1414
<< metal3 >>
rect 655 6580 721 6589
rect 655 6524 660 6580
rect 716 6524 721 6580
rect 354 6202 420 6211
rect 354 6146 359 6202
rect 415 6146 420 6202
rect 354 5446 420 6146
rect 354 5390 359 5446
rect 415 5390 420 5446
rect 354 1414 420 5390
rect 483 5068 549 5077
rect 483 5012 488 5068
rect 544 5012 549 5068
rect 483 4312 549 5012
rect 483 4256 488 4312
rect 544 4256 549 4312
rect 483 3871 549 4256
rect 483 3815 488 3871
rect 544 3815 549 3871
rect 483 3115 549 3815
rect 655 3304 721 6524
rect 655 3248 660 3304
rect 716 3248 721 3304
rect 655 3239 721 3248
rect 827 6580 893 6589
rect 827 6524 832 6580
rect 888 6524 893 6580
rect 827 3304 893 6524
rect 1128 6202 1194 6211
rect 1128 6146 1133 6202
rect 1189 6146 1194 6202
rect 1128 5446 1194 6146
rect 1128 5390 1133 5446
rect 1189 5390 1194 5446
rect 827 3248 832 3304
rect 888 3248 893 3304
rect 827 3239 893 3248
rect 999 5068 1065 5077
rect 999 5012 1004 5068
rect 1060 5012 1065 5068
rect 999 4312 1065 5012
rect 999 4256 1004 4312
rect 1060 4256 1065 4312
rect 999 3493 1065 4256
rect 999 3437 1004 3493
rect 1060 3437 1065 3493
rect 483 3059 488 3115
rect 544 3059 549 3115
rect 483 3050 549 3059
rect 999 3115 1065 3437
rect 999 3059 1004 3115
rect 1060 3059 1065 3115
rect 999 3050 1065 3059
rect 354 1358 359 1414
rect 415 1358 420 1414
rect 354 1349 420 1358
rect 1128 1414 1194 5390
rect 1128 1358 1133 1414
rect 1189 1358 1194 1414
rect 1128 1349 1194 1358
<< labels >>
flabel metal2 s 398 476 1150 532 0 FreeSans 560 0 0 0 VSS
port 1 nsew
flabel metal2 s 398 7658 1150 7714 0 FreeSans 560 0 0 0 VDD
port 2 nsew
flabel metal2 s 484 1358 1064 1414 0 FreeSans 560 0 0 0 clk
port 3 nsew
flabel metal2 s 484 2492 1064 2548 0 FreeSans 560 0 0 0 inn
port 4 nsew
flabel metal2 s 484 2681 1064 2737 0 FreeSans 560 0 0 0 inp
port 5 nsew
flabel metal3 s 999 3050 1065 5077 0 FreeSans 660 90 0 0 outn
port 6 nsew
flabel metal3 s 483 3050 549 5077 0 FreeSans 660 90 0 0 outp
port 7 nsew
flabel metal3 s 655 3239 721 6589 0 FreeSans 660 90 0 0 midn
port 8 nsew
flabel metal3 s 827 3239 893 6589 0 FreeSans 660 90 0 0 midp
port 9 nsew
<< end >>
