magic
tech sky130A
magscale 1 2
timestamp 1645319819
<< checkpaint >>
rect -1000 1662 1609 1713
rect -1318 -1186 1609 1662
rect -1318 -1213 1260 -1186
<< dnwell >>
rect 0 0 260 411
<< pwell >>
rect 0 80 260 362
<< psubdiff >>
rect 0 201 260 336
rect 0 167 79 201
rect 113 167 147 201
rect 181 167 260 201
rect 0 142 260 167
rect 17 108 243 142
rect 0 106 260 108
<< psubdiffcont >>
rect 79 167 113 201
rect 147 167 181 201
rect 0 108 17 142
rect 243 108 260 142
<< poly >>
rect 0 24 260 54
<< locali >>
rect 0 341 70 375
rect 104 341 260 375
rect 0 303 260 341
rect 0 269 70 303
rect 104 269 260 303
rect 0 235 260 269
rect 0 167 79 201
rect 113 167 147 201
rect 181 167 260 201
rect 0 162 260 167
rect 0 142 158 162
rect 17 128 158 142
rect 192 142 260 162
rect 192 128 243 142
rect 17 108 243 128
rect 0 90 260 108
rect 0 56 158 90
rect 192 56 260 90
rect 0 55 260 56
rect 27 3 240 55
<< viali >>
rect 70 341 104 375
rect 70 269 104 303
rect 158 128 192 162
rect 158 56 192 90
<< metal1 >>
rect 0 391 30 411
rect 26 364 30 391
rect 25 340 30 364
rect 0 337 30 340
rect 0 204 18 337
tri 18 325 30 337 nw
rect 62 375 110 411
rect 62 341 70 375
rect 104 341 110 375
tri 50 311 62 323 se
rect 62 311 110 341
rect 50 303 110 311
rect 50 289 70 303
rect 104 289 110 303
rect 50 239 55 289
rect 105 239 110 289
rect 50 231 110 239
tri 18 204 34 220 sw
tri 50 219 62 231 ne
rect 0 146 34 204
rect 0 0 14 146
tri 14 126 34 146 nw
tri 42 76 62 96 se
rect 62 76 110 231
rect 42 34 110 76
rect 42 0 76 34
tri 76 0 110 34 nw
rect 150 311 198 411
rect 230 391 260 411
rect 230 364 234 391
rect 230 340 235 364
rect 230 337 260 340
tri 230 325 242 337 ne
tri 198 311 210 323 sw
rect 150 231 210 311
rect 150 162 198 231
tri 198 219 210 231 nw
rect 150 128 158 162
rect 192 128 198 162
rect 150 90 198 128
tri 226 205 242 221 se
rect 242 205 260 337
rect 226 146 260 205
tri 226 126 246 146 ne
rect 150 56 158 90
rect 192 78 198 90
tri 198 78 216 96 sw
rect 211 76 216 78
tri 216 76 218 78 sw
rect 150 34 161 56
tri 150 28 156 34 ne
rect 156 28 161 34
rect 211 28 218 76
tri 156 0 184 28 ne
rect 184 0 218 28
rect 246 0 260 146
<< via1 >>
rect 0 364 26 391
rect 0 340 25 364
rect 55 269 70 289
rect 70 269 104 289
rect 104 269 105 289
rect 55 239 105 269
rect 234 364 260 391
rect 235 340 260 364
rect 161 56 192 78
rect 192 56 211 78
rect 161 28 211 56
<< metal2 >>
rect 0 391 260 411
rect 26 364 234 391
rect 25 340 235 364
rect 0 320 260 340
rect 0 289 260 292
rect 0 239 55 289
rect 105 239 260 289
rect 0 236 260 239
rect 0 116 260 206
rect 0 78 260 81
rect 0 28 161 78
rect 211 28 260 78
rect 0 4 260 28
<< labels >>
rlabel metal1 s 0 0 14 19 4 VGND
rlabel metal1 s 154 162 198 198 4 VPB
rlabel metal1 s 62 162 106 198 4 VNB
rlabel metal1 s 246 0 260 19 4 VGND
<< end >>
