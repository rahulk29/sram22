.subckt sram_sp_rowtapend_replica VSS VNB
X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 w=0.42 l=0.15
.ends
