magic
tech sky130A
magscale 1 2
timestamp 1644720859
<< checkpaint >>
rect -1020 1461 1597 1733
rect -1290 -1117 1597 1461
rect -1120 -1181 1597 -1117
rect -1120 -1290 1492 -1181
<< dnwell >>
rect 0 0 240 411
<< nwell >>
rect 0 0 96 411
<< pwell >>
rect 114 80 240 362
rect 148 0 228 80
<< nmos >>
rect 174 24 202 52
<< ndiff >>
rect 174 15 202 24
<< ndiffc >>
rect 174 0 202 15
<< psubdiff >>
rect 140 142 240 336
rect 140 108 155 142
rect 189 108 223 142
rect 140 106 240 108
<< nsubdiff >>
rect 0 368 66 375
rect 0 334 17 368
rect 51 334 66 368
rect 0 300 66 334
rect 0 266 17 300
rect 51 266 66 300
rect 0 232 66 266
rect 0 198 17 232
rect 51 198 66 232
rect 0 94 66 198
<< psubdiffcont >>
rect 155 108 189 142
rect 223 108 240 142
<< nsubdiffcont >>
rect 17 334 51 368
rect 17 266 51 300
rect 17 198 51 232
<< poly >>
rect 0 52 240 54
rect 0 24 174 52
rect 202 24 240 52
<< locali >>
rect 0 368 240 375
rect 0 334 17 368
rect 51 334 240 368
rect 0 300 240 334
rect 0 266 17 300
rect 51 266 240 300
rect 0 235 240 266
rect 0 232 68 235
rect 0 198 17 232
rect 51 198 68 232
rect 104 162 240 201
rect 0 142 240 162
rect 0 108 155 142
rect 189 108 223 142
rect 0 55 240 108
rect 14 0 67 15
rect 101 0 174 15
rect 202 0 226 15
<< viali >>
rect 67 0 101 17
<< metal1 >>
rect 0 205 18 411
rect 61 318 97 411
tri 61 310 69 318 ne
tri 18 205 34 221 sw
rect 0 200 34 205
rect 25 150 34 200
rect 0 146 34 150
rect 0 0 14 146
tri 14 126 34 146 nw
rect 69 29 97 318
rect 142 319 178 411
rect 60 17 108 29
rect 60 0 67 17
rect 101 0 108 17
rect 142 0 170 319
tri 170 311 178 319 nw
rect 210 391 240 411
rect 210 364 214 391
rect 210 340 215 364
rect 210 319 240 340
tri 210 303 226 319 ne
rect 226 0 240 319
<< via1 >>
rect 0 150 25 200
rect 214 364 240 391
rect 215 340 240 364
<< metal2 >>
rect 0 391 240 411
rect 0 364 214 391
rect 0 340 215 364
rect 0 320 240 340
rect 0 236 240 292
rect 0 200 240 206
rect 25 150 240 200
rect 0 116 240 150
rect 0 4 240 81
<< labels >>
rlabel metal1 s 69 55 97 81 4 BL1
port 1 se
rlabel metal1 s 0 0 14 19 4 VPWR
port 3 se
rlabel metal1 s 226 0 240 19 4 VGND
port 2 se
rlabel metal1 s 142 55 170 81 4 BL0
port 0 se
<< end >>
