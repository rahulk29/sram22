magic
tech sky130A
timestamp 1643335051
<< nwell >>
rect -47 137 174 300
<< pwell >>
rect -42 0 169 108
<< nmos >>
rect 0 13 15 95
rect 112 13 127 95
<< pmos >>
rect 0 155 15 282
rect 112 155 127 282
<< ndiff >>
rect -29 72 0 95
rect -29 55 -23 72
rect -6 55 0 72
rect -29 38 0 55
rect -29 21 -23 38
rect -6 21 0 38
rect -29 13 0 21
rect 15 74 44 95
rect 15 57 21 74
rect 38 57 44 74
rect 15 40 44 57
rect 15 23 21 40
rect 38 23 44 40
rect 15 13 44 23
rect 83 72 112 95
rect 83 55 89 72
rect 106 55 112 72
rect 83 38 112 55
rect 83 21 89 38
rect 106 21 112 38
rect 83 13 112 21
rect 127 74 156 95
rect 127 57 133 74
rect 150 57 156 74
rect 127 40 156 57
rect 127 23 133 40
rect 150 23 156 40
rect 127 13 156 23
<< pdiff >>
rect -29 248 0 282
rect -29 231 -23 248
rect -6 231 0 248
rect -29 214 0 231
rect -29 197 -23 214
rect -6 197 0 214
rect -29 180 0 197
rect -29 163 -23 180
rect -6 163 0 180
rect -29 155 0 163
rect 15 248 44 282
rect 15 231 21 248
rect 38 231 44 248
rect 15 214 44 231
rect 15 197 21 214
rect 38 197 44 214
rect 15 180 44 197
rect 15 163 21 180
rect 38 163 44 180
rect 15 155 44 163
rect 83 248 112 282
rect 83 231 89 248
rect 106 231 112 248
rect 83 214 112 231
rect 83 197 89 214
rect 106 197 112 214
rect 83 180 112 197
rect 83 163 89 180
rect 106 163 112 180
rect 83 155 112 163
rect 127 248 156 282
rect 127 231 133 248
rect 150 231 156 248
rect 127 214 156 231
rect 127 197 133 214
rect 150 197 156 214
rect 127 180 156 197
rect 127 163 133 180
rect 150 163 156 180
rect 127 155 156 163
<< ndiffc >>
rect -23 55 -6 72
rect -23 21 -6 38
rect 21 57 38 74
rect 21 23 38 40
rect 89 55 106 72
rect 89 21 106 38
rect 133 57 150 74
rect 133 23 150 40
<< pdiffc >>
rect -23 231 -6 248
rect -23 197 -6 214
rect -23 163 -6 180
rect 21 231 38 248
rect 21 197 38 214
rect 21 163 38 180
rect 89 231 106 248
rect 89 197 106 214
rect 89 163 106 180
rect 133 231 150 248
rect 133 197 150 214
rect 133 163 150 180
<< poly >>
rect 0 282 15 295
rect 112 282 127 295
rect 0 139 15 155
rect 112 139 127 155
rect -27 131 15 139
rect -27 114 -22 131
rect -5 114 15 131
rect -27 106 15 114
rect 85 131 127 139
rect 85 114 90 131
rect 107 114 127 131
rect 85 106 127 114
rect 0 95 15 106
rect 112 95 127 106
rect 0 0 15 13
rect 112 0 127 13
<< polycont >>
rect -22 114 -5 131
rect 90 114 107 131
<< locali >>
rect -47 297 174 314
rect -23 248 -6 297
rect -23 214 -6 231
rect -23 180 -6 197
rect -23 155 -6 163
rect 21 248 38 280
rect 21 214 38 231
rect 21 180 38 197
rect -57 114 -22 131
rect -5 114 3 131
rect -57 108 -40 114
rect 21 108 38 163
rect 89 248 106 297
rect 89 214 106 231
rect 89 180 106 197
rect 55 154 72 157
rect 89 155 106 163
rect 133 248 150 280
rect 133 214 150 231
rect 133 180 150 197
rect 55 131 72 137
rect 133 154 150 163
rect 55 114 90 131
rect 107 114 115 131
rect -57 88 -40 91
rect -23 72 -6 95
rect -23 38 -6 55
rect -23 -2 -6 21
rect 21 74 38 91
rect 21 40 38 57
rect 21 15 38 23
rect 89 72 106 95
rect 89 38 106 55
rect 89 -2 106 21
rect 133 74 150 137
rect 133 40 150 57
rect 133 15 150 23
rect -47 -19 174 -2
<< viali >>
rect -57 91 -40 108
rect 55 137 72 154
rect 133 137 150 154
rect 21 91 38 108
<< metal1 >>
rect -83 154 84 157
rect -83 137 55 154
rect 72 137 84 154
rect -83 134 84 137
rect 119 154 174 157
rect 119 137 133 154
rect 150 137 174 154
rect 119 134 174 137
rect -83 108 -28 111
rect -83 91 -57 108
rect -40 91 -28 108
rect -83 88 -28 91
rect 7 108 174 111
rect 7 91 21 108
rect 38 91 174 108
rect 7 88 174 91
<< end >>
