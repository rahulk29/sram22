magic
tech sky130A
magscale 1 2
timestamp 1648174121
<< nwell >>
rect 0 3463 960 7737
<< pwell >>
rect 84 3032 360 3420
rect 600 3032 876 3420
rect 84 1806 360 2194
rect 600 1806 876 2194
rect 84 1332 360 1720
rect 600 1332 876 1720
rect 62 0 898 452
<< nmos >>
rect 164 3058 194 3394
rect 250 3058 280 3394
rect 680 3058 710 3394
rect 766 3058 796 3394
rect 164 1832 194 2168
rect 250 1832 280 2168
rect 680 1832 710 2168
rect 766 1832 796 2168
rect 164 1358 194 1694
rect 250 1358 280 1694
rect 680 1358 710 1694
rect 766 1358 796 1694
<< pmos >>
rect 164 6334 194 6534
rect 250 6334 280 6534
rect 680 6334 710 6534
rect 766 6334 796 6534
rect 164 4892 194 5092
rect 250 4892 280 5092
rect 680 4892 710 5092
rect 766 4892 796 5092
rect 164 3532 194 3932
rect 250 3532 280 3932
rect 680 3532 710 3932
rect 766 3532 796 3932
<< ndiff >>
rect 110 3379 164 3394
rect 110 3345 119 3379
rect 153 3345 164 3379
rect 110 3311 164 3345
rect 110 3277 119 3311
rect 153 3277 164 3311
rect 110 3243 164 3277
rect 110 3209 119 3243
rect 153 3209 164 3243
rect 110 3175 164 3209
rect 110 3141 119 3175
rect 153 3141 164 3175
rect 110 3107 164 3141
rect 110 3073 119 3107
rect 153 3073 164 3107
rect 110 3058 164 3073
rect 194 3379 250 3394
rect 194 3345 205 3379
rect 239 3345 250 3379
rect 194 3311 250 3345
rect 194 3277 205 3311
rect 239 3277 250 3311
rect 194 3243 250 3277
rect 194 3209 205 3243
rect 239 3209 250 3243
rect 194 3175 250 3209
rect 194 3141 205 3175
rect 239 3141 250 3175
rect 194 3107 250 3141
rect 194 3073 205 3107
rect 239 3073 250 3107
rect 194 3058 250 3073
rect 280 3379 334 3394
rect 280 3345 291 3379
rect 325 3345 334 3379
rect 280 3311 334 3345
rect 280 3277 291 3311
rect 325 3277 334 3311
rect 280 3243 334 3277
rect 280 3209 291 3243
rect 325 3209 334 3243
rect 280 3175 334 3209
rect 280 3141 291 3175
rect 325 3141 334 3175
rect 280 3107 334 3141
rect 280 3073 291 3107
rect 325 3073 334 3107
rect 280 3058 334 3073
rect 626 3379 680 3394
rect 626 3345 635 3379
rect 669 3345 680 3379
rect 626 3311 680 3345
rect 626 3277 635 3311
rect 669 3277 680 3311
rect 626 3243 680 3277
rect 626 3209 635 3243
rect 669 3209 680 3243
rect 626 3175 680 3209
rect 626 3141 635 3175
rect 669 3141 680 3175
rect 626 3107 680 3141
rect 626 3073 635 3107
rect 669 3073 680 3107
rect 626 3058 680 3073
rect 710 3379 766 3394
rect 710 3345 721 3379
rect 755 3345 766 3379
rect 710 3311 766 3345
rect 710 3277 721 3311
rect 755 3277 766 3311
rect 710 3243 766 3277
rect 710 3209 721 3243
rect 755 3209 766 3243
rect 710 3175 766 3209
rect 710 3141 721 3175
rect 755 3141 766 3175
rect 710 3107 766 3141
rect 710 3073 721 3107
rect 755 3073 766 3107
rect 710 3058 766 3073
rect 796 3379 850 3394
rect 796 3345 807 3379
rect 841 3345 850 3379
rect 796 3311 850 3345
rect 796 3277 807 3311
rect 841 3277 850 3311
rect 796 3243 850 3277
rect 796 3209 807 3243
rect 841 3209 850 3243
rect 796 3175 850 3209
rect 796 3141 807 3175
rect 841 3141 850 3175
rect 796 3107 850 3141
rect 796 3073 807 3107
rect 841 3073 850 3107
rect 796 3058 850 3073
rect 110 2153 164 2168
rect 110 2119 119 2153
rect 153 2119 164 2153
rect 110 2085 164 2119
rect 110 2051 119 2085
rect 153 2051 164 2085
rect 110 2017 164 2051
rect 110 1983 119 2017
rect 153 1983 164 2017
rect 110 1949 164 1983
rect 110 1915 119 1949
rect 153 1915 164 1949
rect 110 1881 164 1915
rect 110 1847 119 1881
rect 153 1847 164 1881
rect 110 1832 164 1847
rect 194 2153 250 2168
rect 194 2119 205 2153
rect 239 2119 250 2153
rect 194 2085 250 2119
rect 194 2051 205 2085
rect 239 2051 250 2085
rect 194 2017 250 2051
rect 194 1983 205 2017
rect 239 1983 250 2017
rect 194 1949 250 1983
rect 194 1915 205 1949
rect 239 1915 250 1949
rect 194 1881 250 1915
rect 194 1847 205 1881
rect 239 1847 250 1881
rect 194 1832 250 1847
rect 280 2153 334 2168
rect 280 2119 291 2153
rect 325 2119 334 2153
rect 280 2085 334 2119
rect 280 2051 291 2085
rect 325 2051 334 2085
rect 280 2017 334 2051
rect 280 1983 291 2017
rect 325 1983 334 2017
rect 280 1949 334 1983
rect 280 1915 291 1949
rect 325 1915 334 1949
rect 280 1881 334 1915
rect 280 1847 291 1881
rect 325 1847 334 1881
rect 280 1832 334 1847
rect 626 2153 680 2168
rect 626 2119 635 2153
rect 669 2119 680 2153
rect 626 2085 680 2119
rect 626 2051 635 2085
rect 669 2051 680 2085
rect 626 2017 680 2051
rect 626 1983 635 2017
rect 669 1983 680 2017
rect 626 1949 680 1983
rect 626 1915 635 1949
rect 669 1915 680 1949
rect 626 1881 680 1915
rect 626 1847 635 1881
rect 669 1847 680 1881
rect 626 1832 680 1847
rect 710 2153 766 2168
rect 710 2119 721 2153
rect 755 2119 766 2153
rect 710 2085 766 2119
rect 710 2051 721 2085
rect 755 2051 766 2085
rect 710 2017 766 2051
rect 710 1983 721 2017
rect 755 1983 766 2017
rect 710 1949 766 1983
rect 710 1915 721 1949
rect 755 1915 766 1949
rect 710 1881 766 1915
rect 710 1847 721 1881
rect 755 1847 766 1881
rect 710 1832 766 1847
rect 796 2153 850 2168
rect 796 2119 807 2153
rect 841 2119 850 2153
rect 796 2085 850 2119
rect 796 2051 807 2085
rect 841 2051 850 2085
rect 796 2017 850 2051
rect 796 1983 807 2017
rect 841 1983 850 2017
rect 796 1949 850 1983
rect 796 1915 807 1949
rect 841 1915 850 1949
rect 796 1881 850 1915
rect 796 1847 807 1881
rect 841 1847 850 1881
rect 796 1832 850 1847
rect 110 1679 164 1694
rect 110 1645 119 1679
rect 153 1645 164 1679
rect 110 1611 164 1645
rect 110 1577 119 1611
rect 153 1577 164 1611
rect 110 1543 164 1577
rect 110 1509 119 1543
rect 153 1509 164 1543
rect 110 1475 164 1509
rect 110 1441 119 1475
rect 153 1441 164 1475
rect 110 1407 164 1441
rect 110 1373 119 1407
rect 153 1373 164 1407
rect 110 1358 164 1373
rect 194 1679 250 1694
rect 194 1645 205 1679
rect 239 1645 250 1679
rect 194 1611 250 1645
rect 194 1577 205 1611
rect 239 1577 250 1611
rect 194 1543 250 1577
rect 194 1509 205 1543
rect 239 1509 250 1543
rect 194 1475 250 1509
rect 194 1441 205 1475
rect 239 1441 250 1475
rect 194 1407 250 1441
rect 194 1373 205 1407
rect 239 1373 250 1407
rect 194 1358 250 1373
rect 280 1679 334 1694
rect 280 1645 291 1679
rect 325 1645 334 1679
rect 280 1611 334 1645
rect 280 1577 291 1611
rect 325 1577 334 1611
rect 280 1543 334 1577
rect 280 1509 291 1543
rect 325 1509 334 1543
rect 280 1475 334 1509
rect 280 1441 291 1475
rect 325 1441 334 1475
rect 280 1407 334 1441
rect 280 1373 291 1407
rect 325 1373 334 1407
rect 280 1358 334 1373
rect 626 1679 680 1694
rect 626 1645 635 1679
rect 669 1645 680 1679
rect 626 1611 680 1645
rect 626 1577 635 1611
rect 669 1577 680 1611
rect 626 1543 680 1577
rect 626 1509 635 1543
rect 669 1509 680 1543
rect 626 1475 680 1509
rect 626 1441 635 1475
rect 669 1441 680 1475
rect 626 1407 680 1441
rect 626 1373 635 1407
rect 669 1373 680 1407
rect 626 1358 680 1373
rect 710 1679 766 1694
rect 710 1645 721 1679
rect 755 1645 766 1679
rect 710 1611 766 1645
rect 710 1577 721 1611
rect 755 1577 766 1611
rect 710 1543 766 1577
rect 710 1509 721 1543
rect 755 1509 766 1543
rect 710 1475 766 1509
rect 710 1441 721 1475
rect 755 1441 766 1475
rect 710 1407 766 1441
rect 710 1373 721 1407
rect 755 1373 766 1407
rect 710 1358 766 1373
rect 796 1679 850 1694
rect 796 1645 807 1679
rect 841 1645 850 1679
rect 796 1611 850 1645
rect 796 1577 807 1611
rect 841 1577 850 1611
rect 796 1543 850 1577
rect 796 1509 807 1543
rect 841 1509 850 1543
rect 796 1475 850 1509
rect 796 1441 807 1475
rect 841 1441 850 1475
rect 796 1407 850 1441
rect 796 1373 807 1407
rect 841 1373 850 1407
rect 796 1358 850 1373
<< pdiff >>
rect 110 6519 164 6534
rect 110 6485 119 6519
rect 153 6485 164 6519
rect 110 6451 164 6485
rect 110 6417 119 6451
rect 153 6417 164 6451
rect 110 6383 164 6417
rect 110 6349 119 6383
rect 153 6349 164 6383
rect 110 6334 164 6349
rect 194 6519 250 6534
rect 194 6485 205 6519
rect 239 6485 250 6519
rect 194 6451 250 6485
rect 194 6417 205 6451
rect 239 6417 250 6451
rect 194 6383 250 6417
rect 194 6349 205 6383
rect 239 6349 250 6383
rect 194 6334 250 6349
rect 280 6519 334 6534
rect 280 6485 291 6519
rect 325 6485 334 6519
rect 280 6451 334 6485
rect 280 6417 291 6451
rect 325 6417 334 6451
rect 280 6383 334 6417
rect 280 6349 291 6383
rect 325 6349 334 6383
rect 280 6334 334 6349
rect 626 6519 680 6534
rect 626 6485 635 6519
rect 669 6485 680 6519
rect 626 6451 680 6485
rect 626 6417 635 6451
rect 669 6417 680 6451
rect 626 6383 680 6417
rect 626 6349 635 6383
rect 669 6349 680 6383
rect 626 6334 680 6349
rect 710 6519 766 6534
rect 710 6485 721 6519
rect 755 6485 766 6519
rect 710 6451 766 6485
rect 710 6417 721 6451
rect 755 6417 766 6451
rect 710 6383 766 6417
rect 710 6349 721 6383
rect 755 6349 766 6383
rect 710 6334 766 6349
rect 796 6519 850 6534
rect 796 6485 807 6519
rect 841 6485 850 6519
rect 796 6451 850 6485
rect 796 6417 807 6451
rect 841 6417 850 6451
rect 796 6383 850 6417
rect 796 6349 807 6383
rect 841 6349 850 6383
rect 796 6334 850 6349
rect 110 5077 164 5092
rect 110 5043 119 5077
rect 153 5043 164 5077
rect 110 5009 164 5043
rect 110 4975 119 5009
rect 153 4975 164 5009
rect 110 4941 164 4975
rect 110 4907 119 4941
rect 153 4907 164 4941
rect 110 4892 164 4907
rect 194 5077 250 5092
rect 194 5043 205 5077
rect 239 5043 250 5077
rect 194 5009 250 5043
rect 194 4975 205 5009
rect 239 4975 250 5009
rect 194 4941 250 4975
rect 194 4907 205 4941
rect 239 4907 250 4941
rect 194 4892 250 4907
rect 280 5077 334 5092
rect 280 5043 291 5077
rect 325 5043 334 5077
rect 280 5009 334 5043
rect 280 4975 291 5009
rect 325 4975 334 5009
rect 280 4941 334 4975
rect 280 4907 291 4941
rect 325 4907 334 4941
rect 280 4892 334 4907
rect 626 5077 680 5092
rect 626 5043 635 5077
rect 669 5043 680 5077
rect 626 5009 680 5043
rect 626 4975 635 5009
rect 669 4975 680 5009
rect 626 4941 680 4975
rect 626 4907 635 4941
rect 669 4907 680 4941
rect 626 4892 680 4907
rect 710 5077 766 5092
rect 710 5043 721 5077
rect 755 5043 766 5077
rect 710 5009 766 5043
rect 710 4975 721 5009
rect 755 4975 766 5009
rect 710 4941 766 4975
rect 710 4907 721 4941
rect 755 4907 766 4941
rect 710 4892 766 4907
rect 796 5077 850 5092
rect 796 5043 807 5077
rect 841 5043 850 5077
rect 796 5009 850 5043
rect 796 4975 807 5009
rect 841 4975 850 5009
rect 796 4941 850 4975
rect 796 4907 807 4941
rect 841 4907 850 4941
rect 796 4892 850 4907
rect 110 3919 164 3932
rect 110 3885 119 3919
rect 153 3885 164 3919
rect 110 3851 164 3885
rect 110 3817 119 3851
rect 153 3817 164 3851
rect 110 3783 164 3817
rect 110 3749 119 3783
rect 153 3749 164 3783
rect 110 3715 164 3749
rect 110 3681 119 3715
rect 153 3681 164 3715
rect 110 3647 164 3681
rect 110 3613 119 3647
rect 153 3613 164 3647
rect 110 3579 164 3613
rect 110 3545 119 3579
rect 153 3545 164 3579
rect 110 3532 164 3545
rect 194 3919 250 3932
rect 194 3885 205 3919
rect 239 3885 250 3919
rect 194 3851 250 3885
rect 194 3817 205 3851
rect 239 3817 250 3851
rect 194 3783 250 3817
rect 194 3749 205 3783
rect 239 3749 250 3783
rect 194 3715 250 3749
rect 194 3681 205 3715
rect 239 3681 250 3715
rect 194 3647 250 3681
rect 194 3613 205 3647
rect 239 3613 250 3647
rect 194 3579 250 3613
rect 194 3545 205 3579
rect 239 3545 250 3579
rect 194 3532 250 3545
rect 280 3919 334 3932
rect 280 3885 291 3919
rect 325 3885 334 3919
rect 280 3851 334 3885
rect 280 3817 291 3851
rect 325 3817 334 3851
rect 280 3783 334 3817
rect 280 3749 291 3783
rect 325 3749 334 3783
rect 280 3715 334 3749
rect 280 3681 291 3715
rect 325 3681 334 3715
rect 280 3647 334 3681
rect 280 3613 291 3647
rect 325 3613 334 3647
rect 280 3579 334 3613
rect 280 3545 291 3579
rect 325 3545 334 3579
rect 280 3532 334 3545
rect 626 3919 680 3932
rect 626 3885 635 3919
rect 669 3885 680 3919
rect 626 3851 680 3885
rect 626 3817 635 3851
rect 669 3817 680 3851
rect 626 3783 680 3817
rect 626 3749 635 3783
rect 669 3749 680 3783
rect 626 3715 680 3749
rect 626 3681 635 3715
rect 669 3681 680 3715
rect 626 3647 680 3681
rect 626 3613 635 3647
rect 669 3613 680 3647
rect 626 3579 680 3613
rect 626 3545 635 3579
rect 669 3545 680 3579
rect 626 3532 680 3545
rect 710 3919 766 3932
rect 710 3885 721 3919
rect 755 3885 766 3919
rect 710 3851 766 3885
rect 710 3817 721 3851
rect 755 3817 766 3851
rect 710 3783 766 3817
rect 710 3749 721 3783
rect 755 3749 766 3783
rect 710 3715 766 3749
rect 710 3681 721 3715
rect 755 3681 766 3715
rect 710 3647 766 3681
rect 710 3613 721 3647
rect 755 3613 766 3647
rect 710 3579 766 3613
rect 710 3545 721 3579
rect 755 3545 766 3579
rect 710 3532 766 3545
rect 796 3919 850 3932
rect 796 3885 807 3919
rect 841 3885 850 3919
rect 796 3851 850 3885
rect 796 3817 807 3851
rect 841 3817 850 3851
rect 796 3783 850 3817
rect 796 3749 807 3783
rect 841 3749 850 3783
rect 796 3715 850 3749
rect 796 3681 807 3715
rect 841 3681 850 3715
rect 796 3647 850 3681
rect 796 3613 807 3647
rect 841 3613 850 3647
rect 796 3579 850 3613
rect 796 3545 807 3579
rect 841 3545 850 3579
rect 796 3532 850 3545
<< ndiffc >>
rect 119 3345 153 3379
rect 119 3277 153 3311
rect 119 3209 153 3243
rect 119 3141 153 3175
rect 119 3073 153 3107
rect 205 3345 239 3379
rect 205 3277 239 3311
rect 205 3209 239 3243
rect 205 3141 239 3175
rect 205 3073 239 3107
rect 291 3345 325 3379
rect 291 3277 325 3311
rect 291 3209 325 3243
rect 291 3141 325 3175
rect 291 3073 325 3107
rect 635 3345 669 3379
rect 635 3277 669 3311
rect 635 3209 669 3243
rect 635 3141 669 3175
rect 635 3073 669 3107
rect 721 3345 755 3379
rect 721 3277 755 3311
rect 721 3209 755 3243
rect 721 3141 755 3175
rect 721 3073 755 3107
rect 807 3345 841 3379
rect 807 3277 841 3311
rect 807 3209 841 3243
rect 807 3141 841 3175
rect 807 3073 841 3107
rect 119 2119 153 2153
rect 119 2051 153 2085
rect 119 1983 153 2017
rect 119 1915 153 1949
rect 119 1847 153 1881
rect 205 2119 239 2153
rect 205 2051 239 2085
rect 205 1983 239 2017
rect 205 1915 239 1949
rect 205 1847 239 1881
rect 291 2119 325 2153
rect 291 2051 325 2085
rect 291 1983 325 2017
rect 291 1915 325 1949
rect 291 1847 325 1881
rect 635 2119 669 2153
rect 635 2051 669 2085
rect 635 1983 669 2017
rect 635 1915 669 1949
rect 635 1847 669 1881
rect 721 2119 755 2153
rect 721 2051 755 2085
rect 721 1983 755 2017
rect 721 1915 755 1949
rect 721 1847 755 1881
rect 807 2119 841 2153
rect 807 2051 841 2085
rect 807 1983 841 2017
rect 807 1915 841 1949
rect 807 1847 841 1881
rect 119 1645 153 1679
rect 119 1577 153 1611
rect 119 1509 153 1543
rect 119 1441 153 1475
rect 119 1373 153 1407
rect 205 1645 239 1679
rect 205 1577 239 1611
rect 205 1509 239 1543
rect 205 1441 239 1475
rect 205 1373 239 1407
rect 291 1645 325 1679
rect 291 1577 325 1611
rect 291 1509 325 1543
rect 291 1441 325 1475
rect 291 1373 325 1407
rect 635 1645 669 1679
rect 635 1577 669 1611
rect 635 1509 669 1543
rect 635 1441 669 1475
rect 635 1373 669 1407
rect 721 1645 755 1679
rect 721 1577 755 1611
rect 721 1509 755 1543
rect 721 1441 755 1475
rect 721 1373 755 1407
rect 807 1645 841 1679
rect 807 1577 841 1611
rect 807 1509 841 1543
rect 807 1441 841 1475
rect 807 1373 841 1407
<< pdiffc >>
rect 119 6485 153 6519
rect 119 6417 153 6451
rect 119 6349 153 6383
rect 205 6485 239 6519
rect 205 6417 239 6451
rect 205 6349 239 6383
rect 291 6485 325 6519
rect 291 6417 325 6451
rect 291 6349 325 6383
rect 635 6485 669 6519
rect 635 6417 669 6451
rect 635 6349 669 6383
rect 721 6485 755 6519
rect 721 6417 755 6451
rect 721 6349 755 6383
rect 807 6485 841 6519
rect 807 6417 841 6451
rect 807 6349 841 6383
rect 119 5043 153 5077
rect 119 4975 153 5009
rect 119 4907 153 4941
rect 205 5043 239 5077
rect 205 4975 239 5009
rect 205 4907 239 4941
rect 291 5043 325 5077
rect 291 4975 325 5009
rect 291 4907 325 4941
rect 635 5043 669 5077
rect 635 4975 669 5009
rect 635 4907 669 4941
rect 721 5043 755 5077
rect 721 4975 755 5009
rect 721 4907 755 4941
rect 807 5043 841 5077
rect 807 4975 841 5009
rect 807 4907 841 4941
rect 119 3885 153 3919
rect 119 3817 153 3851
rect 119 3749 153 3783
rect 119 3681 153 3715
rect 119 3613 153 3647
rect 119 3545 153 3579
rect 205 3885 239 3919
rect 205 3817 239 3851
rect 205 3749 239 3783
rect 205 3681 239 3715
rect 205 3613 239 3647
rect 205 3545 239 3579
rect 291 3885 325 3919
rect 291 3817 325 3851
rect 291 3749 325 3783
rect 291 3681 325 3715
rect 291 3613 325 3647
rect 291 3545 325 3579
rect 635 3885 669 3919
rect 635 3817 669 3851
rect 635 3749 669 3783
rect 635 3681 669 3715
rect 635 3613 669 3647
rect 635 3545 669 3579
rect 721 3885 755 3919
rect 721 3817 755 3851
rect 721 3749 755 3783
rect 721 3681 755 3715
rect 721 3613 755 3647
rect 721 3545 755 3579
rect 807 3885 841 3919
rect 807 3817 841 3851
rect 807 3749 841 3783
rect 807 3681 841 3715
rect 807 3613 841 3647
rect 807 3545 841 3579
<< psubdiff >>
rect 88 413 872 426
rect 88 379 119 413
rect 153 379 205 413
rect 239 379 291 413
rect 325 379 377 413
rect 411 379 463 413
rect 497 379 549 413
rect 583 379 635 413
rect 669 379 721 413
rect 755 379 807 413
rect 841 379 872 413
rect 88 345 872 379
rect 88 311 119 345
rect 153 311 205 345
rect 239 311 291 345
rect 325 311 377 345
rect 411 311 463 345
rect 497 311 549 345
rect 583 311 635 345
rect 669 311 721 345
rect 755 311 807 345
rect 841 311 872 345
rect 88 277 872 311
rect 88 243 119 277
rect 153 243 205 277
rect 239 243 291 277
rect 325 243 377 277
rect 411 243 463 277
rect 497 243 549 277
rect 583 243 635 277
rect 669 243 721 277
rect 755 243 807 277
rect 841 243 872 277
rect 88 209 872 243
rect 88 175 119 209
rect 153 175 205 209
rect 239 175 291 209
rect 325 175 377 209
rect 411 175 463 209
rect 497 175 549 209
rect 583 175 635 209
rect 669 175 721 209
rect 755 175 807 209
rect 841 175 872 209
rect 88 141 872 175
rect 88 107 119 141
rect 153 107 205 141
rect 239 107 291 141
rect 325 107 377 141
rect 411 107 463 141
rect 497 107 549 141
rect 583 107 635 141
rect 669 107 721 141
rect 755 107 807 141
rect 841 107 872 141
rect 88 73 872 107
rect 88 39 119 73
rect 153 39 205 73
rect 239 39 291 73
rect 325 39 377 73
rect 411 39 463 73
rect 497 39 549 73
rect 583 39 635 73
rect 669 39 721 73
rect 755 39 807 73
rect 841 39 872 73
rect 88 26 872 39
<< nsubdiff >>
rect 88 7529 872 7544
rect 88 7495 119 7529
rect 153 7495 205 7529
rect 239 7495 291 7529
rect 325 7495 377 7529
rect 411 7495 463 7529
rect 497 7495 549 7529
rect 583 7495 635 7529
rect 669 7495 721 7529
rect 755 7495 807 7529
rect 841 7495 872 7529
rect 88 7461 872 7495
rect 88 7427 119 7461
rect 153 7427 205 7461
rect 239 7427 291 7461
rect 325 7427 377 7461
rect 411 7427 463 7461
rect 497 7427 549 7461
rect 583 7427 635 7461
rect 669 7427 721 7461
rect 755 7427 807 7461
rect 841 7427 872 7461
rect 88 7393 872 7427
rect 88 7359 119 7393
rect 153 7359 205 7393
rect 239 7359 291 7393
rect 325 7359 377 7393
rect 411 7359 463 7393
rect 497 7359 549 7393
rect 583 7359 635 7393
rect 669 7359 721 7393
rect 755 7359 807 7393
rect 841 7359 872 7393
rect 88 7325 872 7359
rect 88 7291 119 7325
rect 153 7291 205 7325
rect 239 7291 291 7325
rect 325 7291 377 7325
rect 411 7291 463 7325
rect 497 7291 549 7325
rect 583 7291 635 7325
rect 669 7291 721 7325
rect 755 7291 807 7325
rect 841 7291 872 7325
rect 88 7257 872 7291
rect 88 7223 119 7257
rect 153 7223 205 7257
rect 239 7223 291 7257
rect 325 7223 377 7257
rect 411 7223 463 7257
rect 497 7223 549 7257
rect 583 7223 635 7257
rect 669 7223 721 7257
rect 755 7223 807 7257
rect 841 7223 872 7257
rect 88 7208 872 7223
<< psubdiffcont >>
rect 119 379 153 413
rect 205 379 239 413
rect 291 379 325 413
rect 377 379 411 413
rect 463 379 497 413
rect 549 379 583 413
rect 635 379 669 413
rect 721 379 755 413
rect 807 379 841 413
rect 119 311 153 345
rect 205 311 239 345
rect 291 311 325 345
rect 377 311 411 345
rect 463 311 497 345
rect 549 311 583 345
rect 635 311 669 345
rect 721 311 755 345
rect 807 311 841 345
rect 119 243 153 277
rect 205 243 239 277
rect 291 243 325 277
rect 377 243 411 277
rect 463 243 497 277
rect 549 243 583 277
rect 635 243 669 277
rect 721 243 755 277
rect 807 243 841 277
rect 119 175 153 209
rect 205 175 239 209
rect 291 175 325 209
rect 377 175 411 209
rect 463 175 497 209
rect 549 175 583 209
rect 635 175 669 209
rect 721 175 755 209
rect 807 175 841 209
rect 119 107 153 141
rect 205 107 239 141
rect 291 107 325 141
rect 377 107 411 141
rect 463 107 497 141
rect 549 107 583 141
rect 635 107 669 141
rect 721 107 755 141
rect 807 107 841 141
rect 119 39 153 73
rect 205 39 239 73
rect 291 39 325 73
rect 377 39 411 73
rect 463 39 497 73
rect 549 39 583 73
rect 635 39 669 73
rect 721 39 755 73
rect 807 39 841 73
<< nsubdiffcont >>
rect 119 7495 153 7529
rect 205 7495 239 7529
rect 291 7495 325 7529
rect 377 7495 411 7529
rect 463 7495 497 7529
rect 549 7495 583 7529
rect 635 7495 669 7529
rect 721 7495 755 7529
rect 807 7495 841 7529
rect 119 7427 153 7461
rect 205 7427 239 7461
rect 291 7427 325 7461
rect 377 7427 411 7461
rect 463 7427 497 7461
rect 549 7427 583 7461
rect 635 7427 669 7461
rect 721 7427 755 7461
rect 807 7427 841 7461
rect 119 7359 153 7393
rect 205 7359 239 7393
rect 291 7359 325 7393
rect 377 7359 411 7393
rect 463 7359 497 7393
rect 549 7359 583 7393
rect 635 7359 669 7393
rect 721 7359 755 7393
rect 807 7359 841 7393
rect 119 7291 153 7325
rect 205 7291 239 7325
rect 291 7291 325 7325
rect 377 7291 411 7325
rect 463 7291 497 7325
rect 549 7291 583 7325
rect 635 7291 669 7325
rect 721 7291 755 7325
rect 807 7291 841 7325
rect 119 7223 153 7257
rect 205 7223 239 7257
rect 291 7223 325 7257
rect 377 7223 411 7257
rect 463 7223 497 7257
rect 549 7223 583 7257
rect 635 7223 669 7257
rect 721 7223 755 7257
rect 807 7223 841 7257
<< poly >>
rect 164 6534 194 6560
rect 250 6534 280 6560
rect 680 6534 710 6560
rect 766 6534 796 6560
rect 164 6232 194 6334
rect 250 6232 280 6334
rect 164 6214 280 6232
rect 164 6180 205 6214
rect 239 6180 280 6214
rect 164 6162 280 6180
rect 680 6232 710 6334
rect 766 6232 796 6334
rect 680 6214 796 6232
rect 680 6180 721 6214
rect 755 6180 796 6214
rect 680 6162 796 6180
rect 164 5246 280 5264
rect 164 5212 205 5246
rect 239 5212 280 5246
rect 164 5194 280 5212
rect 164 5092 194 5194
rect 250 5092 280 5194
rect 680 5246 796 5264
rect 680 5212 721 5246
rect 755 5212 796 5246
rect 680 5194 796 5212
rect 680 5092 710 5194
rect 766 5092 796 5194
rect 164 4866 194 4892
rect 250 4866 280 4892
rect 680 4866 710 4892
rect 766 4866 796 4892
rect 164 4086 280 4104
rect 164 4052 205 4086
rect 239 4052 280 4086
rect 164 4034 280 4052
rect 164 3932 194 4034
rect 250 3932 280 4034
rect 680 4086 796 4104
rect 680 4052 721 4086
rect 755 4052 796 4086
rect 680 4034 796 4052
rect 680 3932 710 4034
rect 766 3932 796 4034
rect 164 3506 194 3532
rect 250 3506 280 3532
rect 680 3506 710 3532
rect 766 3506 796 3532
rect 164 3394 194 3420
rect 250 3394 280 3420
rect 680 3394 710 3420
rect 766 3394 796 3420
rect 164 2956 194 3058
rect 250 2956 280 3058
rect 164 2938 280 2956
rect 164 2904 205 2938
rect 239 2904 280 2938
rect 164 2886 280 2904
rect 680 2956 710 3058
rect 766 2956 796 3058
rect 680 2938 796 2956
rect 680 2904 721 2938
rect 755 2904 796 2938
rect 680 2886 796 2904
rect 164 2322 280 2340
rect 164 2288 205 2322
rect 239 2288 280 2322
rect 164 2270 280 2288
rect 164 2168 194 2270
rect 250 2168 280 2270
rect 680 2322 796 2340
rect 680 2288 721 2322
rect 755 2288 796 2322
rect 680 2270 796 2288
rect 680 2168 710 2270
rect 766 2168 796 2270
rect 164 1806 194 1832
rect 250 1806 280 1832
rect 680 1806 710 1832
rect 766 1806 796 1832
rect 164 1694 194 1720
rect 250 1694 280 1720
rect 680 1694 710 1720
rect 766 1694 796 1720
rect 164 1256 194 1358
rect 250 1256 280 1358
rect 164 1238 280 1256
rect 164 1204 205 1238
rect 239 1204 280 1238
rect 164 1186 280 1204
rect 680 1256 710 1358
rect 766 1256 796 1358
rect 680 1238 796 1256
rect 680 1204 721 1238
rect 755 1204 796 1238
rect 680 1186 796 1204
<< polycont >>
rect 205 6180 239 6214
rect 721 6180 755 6214
rect 205 5212 239 5246
rect 721 5212 755 5246
rect 205 4052 239 4086
rect 721 4052 755 4086
rect 205 2904 239 2938
rect 721 2904 755 2938
rect 205 2288 239 2322
rect 721 2288 755 2322
rect 205 1204 239 1238
rect 721 1204 755 1238
<< locali >>
rect 119 7537 153 7545
rect 119 7465 153 7495
rect 119 7393 153 7427
rect 119 7325 153 7359
rect 119 7257 153 7287
rect 119 7207 153 7215
rect 205 7537 239 7545
rect 205 7465 239 7495
rect 205 7393 239 7427
rect 205 7325 239 7359
rect 205 7257 239 7287
rect 205 7207 239 7215
rect 291 7537 325 7545
rect 291 7465 325 7495
rect 291 7393 325 7427
rect 291 7325 325 7359
rect 291 7257 325 7287
rect 291 7207 325 7215
rect 377 7537 411 7545
rect 377 7465 411 7495
rect 377 7393 411 7427
rect 377 7325 411 7359
rect 377 7257 411 7287
rect 377 7207 411 7215
rect 463 7537 497 7545
rect 463 7465 497 7495
rect 463 7393 497 7427
rect 463 7325 497 7359
rect 463 7257 497 7287
rect 463 7207 497 7215
rect 549 7537 583 7545
rect 549 7465 583 7495
rect 549 7393 583 7427
rect 549 7325 583 7359
rect 549 7257 583 7287
rect 549 7207 583 7215
rect 635 7537 669 7545
rect 635 7465 669 7495
rect 635 7393 669 7427
rect 635 7325 669 7359
rect 635 7257 669 7287
rect 635 7207 669 7215
rect 721 7537 755 7545
rect 721 7465 755 7495
rect 721 7393 755 7427
rect 721 7325 755 7359
rect 721 7257 755 7287
rect 721 7207 755 7215
rect 807 7537 841 7545
rect 807 7465 841 7495
rect 807 7393 841 7427
rect 807 7325 841 7359
rect 807 7257 841 7287
rect 807 7207 841 7215
rect 119 6523 153 6535
rect 119 6451 153 6485
rect 119 6383 153 6417
rect 119 6333 153 6345
rect 205 6523 239 6535
rect 205 6451 239 6485
rect 205 6383 239 6417
rect 205 6333 239 6345
rect 291 6523 325 6535
rect 291 6451 325 6485
rect 291 6383 325 6417
rect 291 6333 325 6345
rect 635 6523 669 6535
rect 635 6451 669 6485
rect 635 6383 669 6417
rect 635 6333 669 6345
rect 721 6523 755 6535
rect 721 6451 755 6485
rect 721 6383 755 6417
rect 721 6333 755 6345
rect 807 6523 841 6535
rect 807 6451 841 6485
rect 807 6383 841 6417
rect 807 6333 841 6345
rect 188 6180 205 6214
rect 239 6180 256 6214
rect 704 6180 721 6214
rect 755 6180 772 6214
rect 188 5212 205 5246
rect 239 5212 256 5246
rect 704 5212 721 5246
rect 755 5212 772 5246
rect 119 5081 153 5093
rect 119 5009 153 5043
rect 119 4941 153 4975
rect 119 4891 153 4903
rect 205 5081 239 5093
rect 205 5009 239 5043
rect 205 4941 239 4975
rect 205 4891 239 4903
rect 291 5081 325 5093
rect 291 5009 325 5043
rect 291 4941 325 4975
rect 291 4891 325 4903
rect 635 5081 669 5093
rect 635 5009 669 5043
rect 635 4941 669 4975
rect 635 4891 669 4903
rect 721 5081 755 5093
rect 721 5009 755 5043
rect 721 4941 755 4975
rect 721 4891 755 4903
rect 807 5081 841 5093
rect 807 5009 841 5043
rect 807 4941 841 4975
rect 807 4891 841 4903
rect 188 4052 205 4086
rect 239 4052 256 4086
rect 704 4052 721 4086
rect 755 4052 772 4086
rect 119 3919 153 3935
rect 119 3851 153 3859
rect 119 3783 153 3787
rect 119 3677 153 3681
rect 119 3605 153 3613
rect 119 3529 153 3545
rect 205 3919 239 3935
rect 205 3851 239 3859
rect 205 3783 239 3787
rect 205 3677 239 3681
rect 205 3605 239 3613
rect 205 3529 239 3545
rect 291 3919 325 3935
rect 291 3851 325 3859
rect 291 3783 325 3787
rect 291 3677 325 3681
rect 291 3605 325 3613
rect 291 3529 325 3545
rect 635 3919 669 3935
rect 635 3851 669 3859
rect 635 3783 669 3787
rect 635 3677 669 3681
rect 635 3605 669 3613
rect 635 3529 669 3545
rect 721 3919 755 3935
rect 721 3851 755 3859
rect 721 3783 755 3787
rect 721 3677 755 3681
rect 721 3605 755 3613
rect 721 3529 755 3545
rect 807 3919 841 3935
rect 807 3851 841 3859
rect 807 3783 841 3787
rect 807 3677 841 3681
rect 807 3605 841 3613
rect 807 3529 841 3545
rect 119 3387 153 3395
rect 119 3315 153 3345
rect 119 3243 153 3277
rect 119 3175 153 3209
rect 119 3107 153 3137
rect 119 3057 153 3065
rect 205 3387 239 3395
rect 205 3315 239 3345
rect 205 3243 239 3277
rect 205 3175 239 3209
rect 205 3107 239 3137
rect 205 3057 239 3065
rect 291 3387 325 3395
rect 291 3315 325 3345
rect 291 3243 325 3277
rect 291 3175 325 3209
rect 291 3107 325 3137
rect 291 3057 325 3065
rect 635 3387 669 3395
rect 635 3315 669 3345
rect 635 3243 669 3277
rect 635 3175 669 3209
rect 635 3107 669 3137
rect 635 3057 669 3065
rect 721 3387 755 3395
rect 721 3315 755 3345
rect 721 3243 755 3277
rect 721 3175 755 3209
rect 721 3107 755 3137
rect 721 3057 755 3065
rect 807 3387 841 3395
rect 807 3315 841 3345
rect 807 3243 841 3277
rect 807 3175 841 3209
rect 807 3107 841 3137
rect 807 3057 841 3065
rect 188 2904 205 2938
rect 239 2904 256 2938
rect 704 2904 721 2938
rect 755 2904 772 2938
rect 188 2288 205 2322
rect 239 2288 256 2322
rect 704 2288 721 2322
rect 755 2288 772 2322
rect 119 2161 153 2169
rect 119 2089 153 2119
rect 119 2017 153 2051
rect 119 1949 153 1983
rect 119 1881 153 1911
rect 119 1831 153 1839
rect 205 2161 239 2169
rect 205 2089 239 2119
rect 205 2017 239 2051
rect 205 1949 239 1983
rect 205 1881 239 1911
rect 205 1831 239 1839
rect 291 2161 325 2169
rect 291 2089 325 2119
rect 291 2017 325 2051
rect 291 1949 325 1983
rect 291 1881 325 1911
rect 291 1831 325 1839
rect 635 2161 669 2169
rect 635 2089 669 2119
rect 635 2017 669 2051
rect 635 1949 669 1983
rect 635 1881 669 1911
rect 635 1831 669 1839
rect 721 2161 755 2169
rect 721 2089 755 2119
rect 721 2017 755 2051
rect 721 1949 755 1983
rect 721 1881 755 1911
rect 721 1831 755 1839
rect 807 2161 841 2169
rect 807 2089 841 2119
rect 807 2017 841 2051
rect 807 1949 841 1983
rect 807 1881 841 1911
rect 807 1831 841 1839
rect 119 1687 153 1695
rect 119 1615 153 1645
rect 119 1543 153 1577
rect 119 1475 153 1509
rect 119 1407 153 1437
rect 119 1357 153 1365
rect 205 1687 239 1695
rect 205 1615 239 1645
rect 205 1543 239 1577
rect 205 1475 239 1509
rect 205 1407 239 1437
rect 205 1357 239 1365
rect 291 1687 325 1695
rect 291 1615 325 1645
rect 291 1543 325 1577
rect 291 1475 325 1509
rect 291 1407 325 1437
rect 291 1357 325 1365
rect 635 1687 669 1695
rect 635 1615 669 1645
rect 635 1543 669 1577
rect 635 1475 669 1509
rect 635 1407 669 1437
rect 635 1357 669 1365
rect 721 1687 755 1695
rect 721 1615 755 1645
rect 721 1543 755 1577
rect 721 1475 755 1509
rect 721 1407 755 1437
rect 721 1357 755 1365
rect 807 1687 841 1695
rect 807 1615 841 1645
rect 807 1543 841 1577
rect 807 1475 841 1509
rect 807 1407 841 1437
rect 807 1357 841 1365
rect 188 1204 205 1238
rect 239 1204 256 1238
rect 704 1204 721 1238
rect 755 1204 772 1238
rect 119 413 153 429
rect 119 345 153 353
rect 119 277 153 281
rect 119 171 153 175
rect 119 99 153 107
rect 119 23 153 39
rect 205 413 239 429
rect 205 345 239 353
rect 205 277 239 281
rect 205 171 239 175
rect 205 99 239 107
rect 205 23 239 39
rect 291 413 325 429
rect 291 345 325 353
rect 291 277 325 281
rect 291 171 325 175
rect 291 99 325 107
rect 291 23 325 39
rect 377 413 411 429
rect 377 345 411 353
rect 377 277 411 281
rect 377 171 411 175
rect 377 99 411 107
rect 377 23 411 39
rect 463 413 497 429
rect 463 345 497 353
rect 463 277 497 281
rect 463 171 497 175
rect 463 99 497 107
rect 463 23 497 39
rect 549 413 583 429
rect 549 345 583 353
rect 549 277 583 281
rect 549 171 583 175
rect 549 99 583 107
rect 549 23 583 39
rect 635 413 669 429
rect 635 345 669 353
rect 635 277 669 281
rect 635 171 669 175
rect 635 99 669 107
rect 635 23 669 39
rect 721 413 755 429
rect 721 345 755 353
rect 721 277 755 281
rect 721 171 755 175
rect 721 99 755 107
rect 721 23 755 39
rect 807 413 841 429
rect 807 345 841 353
rect 807 277 841 281
rect 807 171 841 175
rect 807 99 841 107
rect 807 23 841 39
<< viali >>
rect 119 7529 153 7537
rect 119 7503 153 7529
rect 119 7461 153 7465
rect 119 7431 153 7461
rect 119 7359 153 7393
rect 119 7291 153 7321
rect 119 7287 153 7291
rect 119 7223 153 7249
rect 119 7215 153 7223
rect 205 7529 239 7537
rect 205 7503 239 7529
rect 205 7461 239 7465
rect 205 7431 239 7461
rect 205 7359 239 7393
rect 205 7291 239 7321
rect 205 7287 239 7291
rect 205 7223 239 7249
rect 205 7215 239 7223
rect 291 7529 325 7537
rect 291 7503 325 7529
rect 291 7461 325 7465
rect 291 7431 325 7461
rect 291 7359 325 7393
rect 291 7291 325 7321
rect 291 7287 325 7291
rect 291 7223 325 7249
rect 291 7215 325 7223
rect 377 7529 411 7537
rect 377 7503 411 7529
rect 377 7461 411 7465
rect 377 7431 411 7461
rect 377 7359 411 7393
rect 377 7291 411 7321
rect 377 7287 411 7291
rect 377 7223 411 7249
rect 377 7215 411 7223
rect 463 7529 497 7537
rect 463 7503 497 7529
rect 463 7461 497 7465
rect 463 7431 497 7461
rect 463 7359 497 7393
rect 463 7291 497 7321
rect 463 7287 497 7291
rect 463 7223 497 7249
rect 463 7215 497 7223
rect 549 7529 583 7537
rect 549 7503 583 7529
rect 549 7461 583 7465
rect 549 7431 583 7461
rect 549 7359 583 7393
rect 549 7291 583 7321
rect 549 7287 583 7291
rect 549 7223 583 7249
rect 549 7215 583 7223
rect 635 7529 669 7537
rect 635 7503 669 7529
rect 635 7461 669 7465
rect 635 7431 669 7461
rect 635 7359 669 7393
rect 635 7291 669 7321
rect 635 7287 669 7291
rect 635 7223 669 7249
rect 635 7215 669 7223
rect 721 7529 755 7537
rect 721 7503 755 7529
rect 721 7461 755 7465
rect 721 7431 755 7461
rect 721 7359 755 7393
rect 721 7291 755 7321
rect 721 7287 755 7291
rect 721 7223 755 7249
rect 721 7215 755 7223
rect 807 7529 841 7537
rect 807 7503 841 7529
rect 807 7461 841 7465
rect 807 7431 841 7461
rect 807 7359 841 7393
rect 807 7291 841 7321
rect 807 7287 841 7291
rect 807 7223 841 7249
rect 807 7215 841 7223
rect 119 6519 153 6523
rect 119 6489 153 6519
rect 119 6417 153 6451
rect 119 6349 153 6379
rect 119 6345 153 6349
rect 205 6519 239 6523
rect 205 6489 239 6519
rect 205 6417 239 6451
rect 205 6349 239 6379
rect 205 6345 239 6349
rect 291 6519 325 6523
rect 291 6489 325 6519
rect 291 6417 325 6451
rect 291 6349 325 6379
rect 291 6345 325 6349
rect 635 6519 669 6523
rect 635 6489 669 6519
rect 635 6417 669 6451
rect 635 6349 669 6379
rect 635 6345 669 6349
rect 721 6519 755 6523
rect 721 6489 755 6519
rect 721 6417 755 6451
rect 721 6349 755 6379
rect 721 6345 755 6349
rect 807 6519 841 6523
rect 807 6489 841 6519
rect 807 6417 841 6451
rect 807 6349 841 6379
rect 807 6345 841 6349
rect 205 6180 239 6214
rect 721 6180 755 6214
rect 205 5212 239 5246
rect 721 5212 755 5246
rect 119 5077 153 5081
rect 119 5047 153 5077
rect 119 4975 153 5009
rect 119 4907 153 4937
rect 119 4903 153 4907
rect 205 5077 239 5081
rect 205 5047 239 5077
rect 205 4975 239 5009
rect 205 4907 239 4937
rect 205 4903 239 4907
rect 291 5077 325 5081
rect 291 5047 325 5077
rect 291 4975 325 5009
rect 291 4907 325 4937
rect 291 4903 325 4907
rect 635 5077 669 5081
rect 635 5047 669 5077
rect 635 4975 669 5009
rect 635 4907 669 4937
rect 635 4903 669 4907
rect 721 5077 755 5081
rect 721 5047 755 5077
rect 721 4975 755 5009
rect 721 4907 755 4937
rect 721 4903 755 4907
rect 807 5077 841 5081
rect 807 5047 841 5077
rect 807 4975 841 5009
rect 807 4907 841 4937
rect 807 4903 841 4907
rect 205 4052 239 4086
rect 721 4052 755 4086
rect 119 3885 153 3893
rect 119 3859 153 3885
rect 119 3817 153 3821
rect 119 3787 153 3817
rect 119 3715 153 3749
rect 119 3647 153 3677
rect 119 3643 153 3647
rect 119 3579 153 3605
rect 119 3571 153 3579
rect 205 3885 239 3893
rect 205 3859 239 3885
rect 205 3817 239 3821
rect 205 3787 239 3817
rect 205 3715 239 3749
rect 205 3647 239 3677
rect 205 3643 239 3647
rect 205 3579 239 3605
rect 205 3571 239 3579
rect 291 3885 325 3893
rect 291 3859 325 3885
rect 291 3817 325 3821
rect 291 3787 325 3817
rect 291 3715 325 3749
rect 291 3647 325 3677
rect 291 3643 325 3647
rect 291 3579 325 3605
rect 291 3571 325 3579
rect 635 3885 669 3893
rect 635 3859 669 3885
rect 635 3817 669 3821
rect 635 3787 669 3817
rect 635 3715 669 3749
rect 635 3647 669 3677
rect 635 3643 669 3647
rect 635 3579 669 3605
rect 635 3571 669 3579
rect 721 3885 755 3893
rect 721 3859 755 3885
rect 721 3817 755 3821
rect 721 3787 755 3817
rect 721 3715 755 3749
rect 721 3647 755 3677
rect 721 3643 755 3647
rect 721 3579 755 3605
rect 721 3571 755 3579
rect 807 3885 841 3893
rect 807 3859 841 3885
rect 807 3817 841 3821
rect 807 3787 841 3817
rect 807 3715 841 3749
rect 807 3647 841 3677
rect 807 3643 841 3647
rect 807 3579 841 3605
rect 807 3571 841 3579
rect 119 3379 153 3387
rect 119 3353 153 3379
rect 119 3311 153 3315
rect 119 3281 153 3311
rect 119 3209 153 3243
rect 119 3141 153 3171
rect 119 3137 153 3141
rect 119 3073 153 3099
rect 119 3065 153 3073
rect 205 3379 239 3387
rect 205 3353 239 3379
rect 205 3311 239 3315
rect 205 3281 239 3311
rect 205 3209 239 3243
rect 205 3141 239 3171
rect 205 3137 239 3141
rect 205 3073 239 3099
rect 205 3065 239 3073
rect 291 3379 325 3387
rect 291 3353 325 3379
rect 291 3311 325 3315
rect 291 3281 325 3311
rect 291 3209 325 3243
rect 291 3141 325 3171
rect 291 3137 325 3141
rect 291 3073 325 3099
rect 291 3065 325 3073
rect 635 3379 669 3387
rect 635 3353 669 3379
rect 635 3311 669 3315
rect 635 3281 669 3311
rect 635 3209 669 3243
rect 635 3141 669 3171
rect 635 3137 669 3141
rect 635 3073 669 3099
rect 635 3065 669 3073
rect 721 3379 755 3387
rect 721 3353 755 3379
rect 721 3311 755 3315
rect 721 3281 755 3311
rect 721 3209 755 3243
rect 721 3141 755 3171
rect 721 3137 755 3141
rect 721 3073 755 3099
rect 721 3065 755 3073
rect 807 3379 841 3387
rect 807 3353 841 3379
rect 807 3311 841 3315
rect 807 3281 841 3311
rect 807 3209 841 3243
rect 807 3141 841 3171
rect 807 3137 841 3141
rect 807 3073 841 3099
rect 807 3065 841 3073
rect 205 2904 239 2938
rect 721 2904 755 2938
rect 205 2288 239 2322
rect 721 2288 755 2322
rect 119 2153 153 2161
rect 119 2127 153 2153
rect 119 2085 153 2089
rect 119 2055 153 2085
rect 119 1983 153 2017
rect 119 1915 153 1945
rect 119 1911 153 1915
rect 119 1847 153 1873
rect 119 1839 153 1847
rect 205 2153 239 2161
rect 205 2127 239 2153
rect 205 2085 239 2089
rect 205 2055 239 2085
rect 205 1983 239 2017
rect 205 1915 239 1945
rect 205 1911 239 1915
rect 205 1847 239 1873
rect 205 1839 239 1847
rect 291 2153 325 2161
rect 291 2127 325 2153
rect 291 2085 325 2089
rect 291 2055 325 2085
rect 291 1983 325 2017
rect 291 1915 325 1945
rect 291 1911 325 1915
rect 291 1847 325 1873
rect 291 1839 325 1847
rect 635 2153 669 2161
rect 635 2127 669 2153
rect 635 2085 669 2089
rect 635 2055 669 2085
rect 635 1983 669 2017
rect 635 1915 669 1945
rect 635 1911 669 1915
rect 635 1847 669 1873
rect 635 1839 669 1847
rect 721 2153 755 2161
rect 721 2127 755 2153
rect 721 2085 755 2089
rect 721 2055 755 2085
rect 721 1983 755 2017
rect 721 1915 755 1945
rect 721 1911 755 1915
rect 721 1847 755 1873
rect 721 1839 755 1847
rect 807 2153 841 2161
rect 807 2127 841 2153
rect 807 2085 841 2089
rect 807 2055 841 2085
rect 807 1983 841 2017
rect 807 1915 841 1945
rect 807 1911 841 1915
rect 807 1847 841 1873
rect 807 1839 841 1847
rect 119 1679 153 1687
rect 119 1653 153 1679
rect 119 1611 153 1615
rect 119 1581 153 1611
rect 119 1509 153 1543
rect 119 1441 153 1471
rect 119 1437 153 1441
rect 119 1373 153 1399
rect 119 1365 153 1373
rect 205 1679 239 1687
rect 205 1653 239 1679
rect 205 1611 239 1615
rect 205 1581 239 1611
rect 205 1509 239 1543
rect 205 1441 239 1471
rect 205 1437 239 1441
rect 205 1373 239 1399
rect 205 1365 239 1373
rect 291 1679 325 1687
rect 291 1653 325 1679
rect 291 1611 325 1615
rect 291 1581 325 1611
rect 291 1509 325 1543
rect 291 1441 325 1471
rect 291 1437 325 1441
rect 291 1373 325 1399
rect 291 1365 325 1373
rect 635 1679 669 1687
rect 635 1653 669 1679
rect 635 1611 669 1615
rect 635 1581 669 1611
rect 635 1509 669 1543
rect 635 1441 669 1471
rect 635 1437 669 1441
rect 635 1373 669 1399
rect 635 1365 669 1373
rect 721 1679 755 1687
rect 721 1653 755 1679
rect 721 1611 755 1615
rect 721 1581 755 1611
rect 721 1509 755 1543
rect 721 1441 755 1471
rect 721 1437 755 1441
rect 721 1373 755 1399
rect 721 1365 755 1373
rect 807 1679 841 1687
rect 807 1653 841 1679
rect 807 1611 841 1615
rect 807 1581 841 1611
rect 807 1509 841 1543
rect 807 1441 841 1471
rect 807 1437 841 1441
rect 807 1373 841 1399
rect 807 1365 841 1373
rect 205 1204 239 1238
rect 721 1204 755 1238
rect 119 379 153 387
rect 119 353 153 379
rect 119 311 153 315
rect 119 281 153 311
rect 119 209 153 243
rect 119 141 153 171
rect 119 137 153 141
rect 119 73 153 99
rect 119 65 153 73
rect 205 379 239 387
rect 205 353 239 379
rect 205 311 239 315
rect 205 281 239 311
rect 205 209 239 243
rect 205 141 239 171
rect 205 137 239 141
rect 205 73 239 99
rect 205 65 239 73
rect 291 379 325 387
rect 291 353 325 379
rect 291 311 325 315
rect 291 281 325 311
rect 291 209 325 243
rect 291 141 325 171
rect 291 137 325 141
rect 291 73 325 99
rect 291 65 325 73
rect 377 379 411 387
rect 377 353 411 379
rect 377 311 411 315
rect 377 281 411 311
rect 377 209 411 243
rect 377 141 411 171
rect 377 137 411 141
rect 377 73 411 99
rect 377 65 411 73
rect 463 379 497 387
rect 463 353 497 379
rect 463 311 497 315
rect 463 281 497 311
rect 463 209 497 243
rect 463 141 497 171
rect 463 137 497 141
rect 463 73 497 99
rect 463 65 497 73
rect 549 379 583 387
rect 549 353 583 379
rect 549 311 583 315
rect 549 281 583 311
rect 549 209 583 243
rect 549 141 583 171
rect 549 137 583 141
rect 549 73 583 99
rect 549 65 583 73
rect 635 379 669 387
rect 635 353 669 379
rect 635 311 669 315
rect 635 281 669 311
rect 635 209 669 243
rect 635 141 669 171
rect 635 137 669 141
rect 635 73 669 99
rect 635 65 669 73
rect 721 379 755 387
rect 721 353 755 379
rect 721 311 755 315
rect 721 281 755 311
rect 721 209 755 243
rect 721 141 755 171
rect 721 137 755 141
rect 721 73 755 99
rect 721 65 755 73
rect 807 379 841 387
rect 807 353 841 379
rect 807 311 841 315
rect 807 281 841 311
rect 807 209 841 243
rect 807 141 841 171
rect 807 137 841 141
rect 807 73 841 99
rect 807 65 841 73
<< metal1 >>
rect 110 7543 162 7549
rect 110 7465 162 7491
rect 110 7431 119 7465
rect 153 7431 162 7465
rect 110 7393 162 7431
rect 110 7359 119 7393
rect 153 7359 162 7393
rect 110 7321 162 7359
rect 110 7287 119 7321
rect 153 7287 162 7321
rect 110 7249 162 7287
rect 110 7215 119 7249
rect 153 7215 162 7249
rect 110 6523 162 7215
rect 196 7543 248 7549
rect 196 7465 248 7491
rect 196 7431 205 7465
rect 239 7431 248 7465
rect 196 7393 248 7431
rect 196 7359 205 7393
rect 239 7359 248 7393
rect 196 7321 248 7359
rect 196 7287 205 7321
rect 239 7287 248 7321
rect 196 7249 248 7287
rect 196 7215 205 7249
rect 239 7215 248 7249
rect 196 7203 248 7215
rect 282 7543 334 7549
rect 282 7465 334 7491
rect 282 7431 291 7465
rect 325 7431 334 7465
rect 282 7393 334 7431
rect 282 7359 291 7393
rect 325 7359 334 7393
rect 282 7321 334 7359
rect 282 7287 291 7321
rect 325 7287 334 7321
rect 282 7249 334 7287
rect 282 7215 291 7249
rect 325 7215 334 7249
rect 110 6489 119 6523
rect 153 6489 162 6523
rect 110 6451 162 6489
rect 110 6417 119 6451
rect 153 6417 162 6451
rect 110 6379 162 6417
rect 110 6345 119 6379
rect 153 6345 162 6379
rect 110 5081 162 6345
rect 196 6523 248 6535
rect 196 6489 205 6523
rect 239 6489 248 6523
rect 196 6451 248 6489
rect 196 6417 205 6451
rect 239 6417 248 6451
rect 196 6409 248 6417
rect 196 6345 205 6357
rect 239 6345 248 6357
rect 196 6333 248 6345
rect 282 6523 334 7215
rect 368 7543 420 7549
rect 368 7465 420 7491
rect 368 7431 377 7465
rect 411 7431 420 7465
rect 368 7393 420 7431
rect 368 7359 377 7393
rect 411 7359 420 7393
rect 368 7321 420 7359
rect 368 7287 377 7321
rect 411 7287 420 7321
rect 368 7249 420 7287
rect 368 7215 377 7249
rect 411 7215 420 7249
rect 368 7203 420 7215
rect 454 7543 506 7549
rect 454 7465 506 7491
rect 454 7431 463 7465
rect 497 7431 506 7465
rect 454 7393 506 7431
rect 454 7359 463 7393
rect 497 7359 506 7393
rect 454 7321 506 7359
rect 454 7287 463 7321
rect 497 7287 506 7321
rect 454 7249 506 7287
rect 454 7215 463 7249
rect 497 7215 506 7249
rect 454 7203 506 7215
rect 540 7543 592 7549
rect 540 7465 592 7491
rect 540 7431 549 7465
rect 583 7431 592 7465
rect 540 7393 592 7431
rect 540 7359 549 7393
rect 583 7359 592 7393
rect 540 7321 592 7359
rect 540 7287 549 7321
rect 583 7287 592 7321
rect 540 7249 592 7287
rect 540 7215 549 7249
rect 583 7215 592 7249
rect 540 7203 592 7215
rect 626 7543 678 7549
rect 626 7465 678 7491
rect 626 7431 635 7465
rect 669 7431 678 7465
rect 626 7393 678 7431
rect 626 7359 635 7393
rect 669 7359 678 7393
rect 626 7321 678 7359
rect 626 7287 635 7321
rect 669 7287 678 7321
rect 626 7249 678 7287
rect 626 7215 635 7249
rect 669 7215 678 7249
rect 392 6986 456 6992
rect 392 6934 398 6986
rect 450 6934 456 6986
rect 392 6928 456 6934
rect 504 6986 568 6992
rect 504 6934 510 6986
rect 562 6934 568 6986
rect 504 6928 568 6934
rect 282 6489 291 6523
rect 325 6489 334 6523
rect 282 6451 334 6489
rect 282 6417 291 6451
rect 325 6417 334 6451
rect 282 6379 334 6417
rect 282 6345 291 6379
rect 325 6345 334 6379
rect 196 6214 248 6226
rect 196 6180 205 6214
rect 239 6180 248 6214
rect 196 6031 248 6180
rect 196 5973 248 5979
rect 196 5275 248 5281
rect 196 5212 205 5223
rect 239 5212 248 5223
rect 196 5200 248 5212
rect 110 5047 119 5081
rect 153 5047 162 5081
rect 110 5009 162 5047
rect 110 4975 119 5009
rect 153 4975 162 5009
rect 110 4937 162 4975
rect 110 4903 119 4937
rect 153 4903 162 4937
rect 110 3893 162 4903
rect 196 5081 248 5093
rect 196 5047 205 5081
rect 239 5047 248 5081
rect 196 5009 248 5047
rect 196 4975 205 5009
rect 239 4975 248 5009
rect 196 4937 248 4975
rect 196 4903 205 4937
rect 239 4903 248 4937
rect 196 4897 248 4903
rect 196 4839 248 4845
rect 282 5081 334 6345
rect 282 5047 291 5081
rect 325 5047 334 5081
rect 282 5009 334 5047
rect 282 4975 291 5009
rect 325 4975 334 5009
rect 282 4937 334 4975
rect 282 4903 291 4937
rect 325 4903 334 4937
rect 196 4141 248 4147
rect 196 4086 248 4089
rect 196 4052 205 4086
rect 239 4052 248 4086
rect 196 4040 248 4052
rect 110 3859 119 3893
rect 153 3859 162 3893
rect 110 3821 162 3859
rect 110 3787 119 3821
rect 153 3787 162 3821
rect 110 3749 162 3787
rect 110 3715 119 3749
rect 153 3715 162 3749
rect 110 3677 162 3715
rect 110 3643 119 3677
rect 153 3643 162 3677
rect 110 3605 162 3643
rect 110 3571 119 3605
rect 153 3571 162 3605
rect 110 3559 162 3571
rect 196 3893 248 3905
rect 196 3859 205 3893
rect 239 3859 248 3893
rect 196 3821 248 3859
rect 196 3787 205 3821
rect 239 3787 248 3821
rect 196 3749 248 3787
rect 196 3715 205 3749
rect 239 3715 248 3749
rect 196 3677 248 3715
rect 196 3643 205 3677
rect 239 3643 248 3677
rect 196 3605 248 3643
rect 196 3571 205 3605
rect 239 3571 248 3605
rect 110 3387 162 3399
rect 110 3353 119 3387
rect 153 3353 162 3387
rect 110 3315 162 3353
rect 110 3281 119 3315
rect 153 3281 162 3315
rect 110 3243 162 3281
rect 110 3209 119 3243
rect 153 3209 162 3243
rect 110 3171 162 3209
rect 110 3137 119 3171
rect 153 3137 162 3171
rect 110 3133 162 3137
rect 110 3065 119 3081
rect 153 3065 162 3081
rect 110 2161 162 3065
rect 196 3387 248 3571
rect 282 3893 334 4903
rect 282 3859 291 3893
rect 325 3859 334 3893
rect 282 3821 334 3859
rect 282 3787 291 3821
rect 325 3787 334 3821
rect 282 3749 334 3787
rect 282 3715 291 3749
rect 325 3715 334 3749
rect 282 3677 334 3715
rect 282 3643 291 3677
rect 325 3643 334 3677
rect 282 3605 334 3643
rect 282 3571 291 3605
rect 325 3571 334 3605
rect 282 3559 334 3571
rect 196 3353 205 3387
rect 239 3353 248 3387
rect 196 3322 248 3353
rect 196 3243 248 3270
rect 196 3209 205 3243
rect 239 3209 248 3243
rect 196 3171 248 3209
rect 196 3137 205 3171
rect 239 3137 248 3171
rect 196 3099 248 3137
rect 196 3065 205 3099
rect 239 3065 248 3099
rect 196 3053 248 3065
rect 282 3387 334 3399
rect 282 3353 291 3387
rect 325 3353 334 3387
rect 282 3315 334 3353
rect 282 3281 291 3315
rect 325 3281 334 3315
rect 282 3243 334 3281
rect 282 3209 291 3243
rect 325 3209 334 3243
rect 282 3171 334 3209
rect 282 3137 291 3171
rect 325 3137 334 3171
rect 282 3133 334 3137
rect 282 3065 291 3081
rect 325 3065 334 3081
rect 196 2944 248 2950
rect 196 2886 248 2892
rect 196 2566 248 2572
rect 196 2322 248 2514
rect 196 2288 205 2322
rect 239 2288 248 2322
rect 196 2276 248 2288
rect 110 2127 119 2161
rect 153 2127 162 2161
rect 110 2089 162 2127
rect 110 2055 119 2089
rect 153 2055 162 2089
rect 110 2017 162 2055
rect 110 1983 119 2017
rect 153 1983 162 2017
rect 110 1945 162 1983
rect 110 1911 119 1945
rect 153 1911 162 1945
rect 110 1873 162 1911
rect 110 1839 119 1873
rect 153 1839 162 1873
rect 110 1827 162 1839
rect 196 2161 248 2173
rect 196 2127 205 2161
rect 239 2127 248 2161
rect 196 2089 248 2127
rect 196 2055 205 2089
rect 239 2055 248 2089
rect 196 2017 248 2055
rect 196 1983 205 2017
rect 239 1983 248 2017
rect 196 1945 248 1983
rect 196 1936 205 1945
rect 239 1936 248 1945
rect 196 1873 248 1884
rect 196 1839 205 1873
rect 239 1839 248 1873
rect 110 1687 162 1699
rect 110 1653 119 1687
rect 153 1653 162 1687
rect 110 1615 162 1653
rect 110 1581 119 1615
rect 153 1581 162 1615
rect 110 1543 162 1581
rect 110 1509 119 1543
rect 153 1509 162 1543
rect 110 1471 162 1509
rect 110 1437 119 1471
rect 153 1437 162 1471
rect 110 1399 162 1437
rect 110 1365 119 1399
rect 153 1365 162 1399
rect 110 387 162 1365
rect 196 1687 248 1839
rect 282 2161 334 3065
rect 398 2566 450 6928
rect 398 2503 450 2514
rect 510 2377 562 6928
rect 626 6523 678 7215
rect 712 7543 764 7549
rect 712 7465 764 7491
rect 712 7431 721 7465
rect 755 7431 764 7465
rect 712 7393 764 7431
rect 712 7359 721 7393
rect 755 7359 764 7393
rect 712 7321 764 7359
rect 712 7287 721 7321
rect 755 7287 764 7321
rect 712 7249 764 7287
rect 712 7215 721 7249
rect 755 7215 764 7249
rect 712 7203 764 7215
rect 798 7543 850 7549
rect 798 7465 850 7491
rect 798 7431 807 7465
rect 841 7431 850 7465
rect 798 7393 850 7431
rect 798 7359 807 7393
rect 841 7359 850 7393
rect 798 7321 850 7359
rect 798 7287 807 7321
rect 841 7287 850 7321
rect 798 7249 850 7287
rect 798 7215 807 7249
rect 841 7215 850 7249
rect 626 6489 635 6523
rect 669 6489 678 6523
rect 626 6451 678 6489
rect 626 6417 635 6451
rect 669 6417 678 6451
rect 626 6379 678 6417
rect 626 6345 635 6379
rect 669 6345 678 6379
rect 626 5081 678 6345
rect 712 6523 764 6535
rect 712 6489 721 6523
rect 755 6489 764 6523
rect 712 6451 764 6489
rect 712 6417 721 6451
rect 755 6417 764 6451
rect 712 6409 764 6417
rect 712 6345 721 6357
rect 755 6345 764 6357
rect 712 6333 764 6345
rect 798 6523 850 7215
rect 798 6489 807 6523
rect 841 6489 850 6523
rect 798 6451 850 6489
rect 798 6417 807 6451
rect 841 6417 850 6451
rect 798 6379 850 6417
rect 798 6345 807 6379
rect 841 6345 850 6379
rect 712 6214 764 6226
rect 712 6180 721 6214
rect 755 6180 764 6214
rect 712 6031 764 6180
rect 712 5973 764 5979
rect 712 5275 764 5281
rect 712 5212 721 5223
rect 755 5212 764 5223
rect 712 5200 764 5212
rect 626 5047 635 5081
rect 669 5047 678 5081
rect 626 5009 678 5047
rect 626 4975 635 5009
rect 669 4975 678 5009
rect 626 4937 678 4975
rect 626 4903 635 4937
rect 669 4903 678 4937
rect 626 3893 678 4903
rect 712 5081 764 5093
rect 712 5047 721 5081
rect 755 5047 764 5081
rect 712 5009 764 5047
rect 712 4975 721 5009
rect 755 4975 764 5009
rect 712 4937 764 4975
rect 712 4903 721 4937
rect 755 4903 764 4937
rect 712 4897 764 4903
rect 712 4839 764 4845
rect 798 5081 850 6345
rect 798 5047 807 5081
rect 841 5047 850 5081
rect 798 5009 850 5047
rect 798 4975 807 5009
rect 841 4975 850 5009
rect 798 4937 850 4975
rect 798 4903 807 4937
rect 841 4903 850 4937
rect 712 4141 764 4147
rect 712 4086 764 4089
rect 712 4052 721 4086
rect 755 4052 764 4086
rect 712 4040 764 4052
rect 626 3859 635 3893
rect 669 3859 678 3893
rect 626 3821 678 3859
rect 626 3787 635 3821
rect 669 3787 678 3821
rect 626 3749 678 3787
rect 626 3715 635 3749
rect 669 3715 678 3749
rect 626 3677 678 3715
rect 626 3643 635 3677
rect 669 3643 678 3677
rect 626 3605 678 3643
rect 626 3571 635 3605
rect 669 3571 678 3605
rect 626 3559 678 3571
rect 712 3893 764 3905
rect 712 3859 721 3893
rect 755 3859 764 3893
rect 712 3821 764 3859
rect 712 3787 721 3821
rect 755 3787 764 3821
rect 712 3749 764 3787
rect 712 3715 721 3749
rect 755 3715 764 3749
rect 712 3700 764 3715
rect 712 3643 721 3648
rect 755 3643 764 3648
rect 712 3605 764 3643
rect 712 3571 721 3605
rect 755 3571 764 3605
rect 510 2315 562 2325
rect 626 3387 678 3399
rect 626 3353 635 3387
rect 669 3353 678 3387
rect 626 3315 678 3353
rect 626 3281 635 3315
rect 669 3281 678 3315
rect 626 3243 678 3281
rect 626 3209 635 3243
rect 669 3209 678 3243
rect 626 3171 678 3209
rect 626 3137 635 3171
rect 669 3137 678 3171
rect 626 3133 678 3137
rect 626 3065 635 3081
rect 669 3065 678 3081
rect 282 2127 291 2161
rect 325 2127 334 2161
rect 282 2089 334 2127
rect 282 2055 291 2089
rect 325 2055 334 2089
rect 282 2017 334 2055
rect 282 1983 291 2017
rect 325 1983 334 2017
rect 282 1945 334 1983
rect 282 1911 291 1945
rect 325 1911 334 1945
rect 282 1873 334 1911
rect 282 1839 291 1873
rect 325 1839 334 1873
rect 282 1827 334 1839
rect 626 2161 678 3065
rect 712 3387 764 3571
rect 798 3893 850 4903
rect 798 3859 807 3893
rect 841 3859 850 3893
rect 798 3821 850 3859
rect 798 3787 807 3821
rect 841 3787 850 3821
rect 798 3749 850 3787
rect 798 3715 807 3749
rect 841 3715 850 3749
rect 798 3677 850 3715
rect 798 3643 807 3677
rect 841 3643 850 3677
rect 798 3605 850 3643
rect 798 3571 807 3605
rect 841 3571 850 3605
rect 798 3559 850 3571
rect 712 3353 721 3387
rect 755 3353 764 3387
rect 712 3315 764 3353
rect 712 3281 721 3315
rect 755 3281 764 3315
rect 712 3243 764 3281
rect 712 3209 721 3243
rect 755 3209 764 3243
rect 712 3171 764 3209
rect 712 3137 721 3171
rect 755 3137 764 3171
rect 712 3099 764 3137
rect 712 3065 721 3099
rect 755 3065 764 3099
rect 712 3053 764 3065
rect 798 3387 850 3399
rect 798 3353 807 3387
rect 841 3353 850 3387
rect 798 3315 850 3353
rect 798 3281 807 3315
rect 841 3281 850 3315
rect 798 3243 850 3281
rect 798 3209 807 3243
rect 841 3209 850 3243
rect 798 3171 850 3209
rect 798 3137 807 3171
rect 841 3137 850 3171
rect 798 3133 850 3137
rect 798 3065 807 3081
rect 841 3065 850 3081
rect 712 2944 764 2950
rect 712 2886 764 2892
rect 712 2377 764 2572
rect 712 2322 764 2325
rect 712 2288 721 2322
rect 755 2288 764 2322
rect 712 2276 764 2288
rect 626 2127 635 2161
rect 669 2127 678 2161
rect 626 2089 678 2127
rect 626 2055 635 2089
rect 669 2055 678 2089
rect 626 2017 678 2055
rect 626 1983 635 2017
rect 669 1983 678 2017
rect 626 1945 678 1983
rect 626 1911 635 1945
rect 669 1911 678 1945
rect 626 1873 678 1911
rect 626 1839 635 1873
rect 669 1839 678 1873
rect 626 1827 678 1839
rect 712 2161 764 2173
rect 712 2127 721 2161
rect 755 2127 764 2161
rect 712 2089 764 2127
rect 712 2055 721 2089
rect 755 2055 764 2089
rect 712 2017 764 2055
rect 712 1983 721 2017
rect 755 1983 764 2017
rect 712 1945 764 1983
rect 712 1936 721 1945
rect 755 1936 764 1945
rect 712 1873 764 1884
rect 712 1839 721 1873
rect 755 1839 764 1873
rect 196 1653 205 1687
rect 239 1653 248 1687
rect 196 1615 248 1653
rect 196 1581 205 1615
rect 239 1581 248 1615
rect 196 1543 248 1581
rect 196 1509 205 1543
rect 239 1509 248 1543
rect 196 1471 248 1509
rect 196 1437 205 1471
rect 239 1437 248 1471
rect 196 1399 248 1437
rect 196 1365 205 1399
rect 239 1365 248 1399
rect 196 1353 248 1365
rect 282 1687 334 1699
rect 282 1653 291 1687
rect 325 1653 334 1687
rect 282 1615 334 1653
rect 282 1581 291 1615
rect 325 1581 334 1615
rect 282 1543 334 1581
rect 282 1509 291 1543
rect 325 1509 334 1543
rect 282 1471 334 1509
rect 282 1437 291 1471
rect 325 1437 334 1471
rect 282 1399 334 1437
rect 282 1365 291 1399
rect 325 1365 334 1399
rect 196 1243 248 1250
rect 196 1185 248 1191
rect 110 361 119 387
rect 153 361 162 387
rect 110 281 119 309
rect 153 281 162 309
rect 110 243 162 281
rect 110 209 119 243
rect 153 209 162 243
rect 110 171 162 209
rect 110 137 119 171
rect 153 137 162 171
rect 110 99 162 137
rect 110 65 119 99
rect 153 65 162 99
rect 110 53 162 65
rect 196 387 248 399
rect 196 361 205 387
rect 239 361 248 387
rect 196 281 205 309
rect 239 281 248 309
rect 196 243 248 281
rect 196 209 205 243
rect 239 209 248 243
rect 196 171 248 209
rect 196 137 205 171
rect 239 137 248 171
rect 196 99 248 137
rect 196 65 205 99
rect 239 65 248 99
rect 196 53 248 65
rect 282 387 334 1365
rect 626 1687 678 1699
rect 626 1653 635 1687
rect 669 1653 678 1687
rect 626 1615 678 1653
rect 626 1581 635 1615
rect 669 1581 678 1615
rect 626 1543 678 1581
rect 626 1509 635 1543
rect 669 1509 678 1543
rect 626 1471 678 1509
rect 626 1437 635 1471
rect 669 1437 678 1471
rect 626 1399 678 1437
rect 626 1365 635 1399
rect 669 1365 678 1399
rect 282 361 291 387
rect 325 361 334 387
rect 282 281 291 309
rect 325 281 334 309
rect 282 243 334 281
rect 282 209 291 243
rect 325 209 334 243
rect 282 171 334 209
rect 282 137 291 171
rect 325 137 334 171
rect 282 99 334 137
rect 282 65 291 99
rect 325 65 334 99
rect 282 53 334 65
rect 368 387 420 399
rect 368 361 377 387
rect 411 361 420 387
rect 368 281 377 309
rect 411 281 420 309
rect 368 243 420 281
rect 368 209 377 243
rect 411 209 420 243
rect 368 171 420 209
rect 368 137 377 171
rect 411 137 420 171
rect 368 99 420 137
rect 368 65 377 99
rect 411 65 420 99
rect 368 53 420 65
rect 454 387 506 399
rect 454 361 463 387
rect 497 361 506 387
rect 454 281 463 309
rect 497 281 506 309
rect 454 243 506 281
rect 454 209 463 243
rect 497 209 506 243
rect 454 171 506 209
rect 454 137 463 171
rect 497 137 506 171
rect 454 99 506 137
rect 454 65 463 99
rect 497 65 506 99
rect 454 53 506 65
rect 540 387 592 399
rect 540 361 549 387
rect 583 361 592 387
rect 540 281 549 309
rect 583 281 592 309
rect 540 243 592 281
rect 540 209 549 243
rect 583 209 592 243
rect 540 171 592 209
rect 540 137 549 171
rect 583 137 592 171
rect 540 99 592 137
rect 540 65 549 99
rect 583 65 592 99
rect 540 53 592 65
rect 626 387 678 1365
rect 712 1687 764 1839
rect 798 2161 850 3065
rect 798 2127 807 2161
rect 841 2127 850 2161
rect 798 2089 850 2127
rect 798 2055 807 2089
rect 841 2055 850 2089
rect 798 2017 850 2055
rect 798 1983 807 2017
rect 841 1983 850 2017
rect 798 1945 850 1983
rect 798 1911 807 1945
rect 841 1911 850 1945
rect 798 1873 850 1911
rect 798 1839 807 1873
rect 841 1839 850 1873
rect 798 1827 850 1839
rect 712 1653 721 1687
rect 755 1653 764 1687
rect 712 1615 764 1653
rect 712 1581 721 1615
rect 755 1581 764 1615
rect 712 1543 764 1581
rect 712 1509 721 1543
rect 755 1509 764 1543
rect 712 1471 764 1509
rect 712 1437 721 1471
rect 755 1437 764 1471
rect 712 1399 764 1437
rect 712 1365 721 1399
rect 755 1365 764 1399
rect 712 1353 764 1365
rect 798 1687 850 1699
rect 798 1653 807 1687
rect 841 1653 850 1687
rect 798 1615 850 1653
rect 798 1581 807 1615
rect 841 1581 850 1615
rect 798 1543 850 1581
rect 798 1509 807 1543
rect 841 1509 850 1543
rect 798 1471 850 1509
rect 798 1437 807 1471
rect 841 1437 850 1471
rect 798 1399 850 1437
rect 798 1365 807 1399
rect 841 1365 850 1399
rect 712 1243 764 1250
rect 712 1185 764 1191
rect 626 361 635 387
rect 669 361 678 387
rect 626 281 635 309
rect 669 281 678 309
rect 626 243 678 281
rect 626 209 635 243
rect 669 209 678 243
rect 626 171 678 209
rect 626 137 635 171
rect 669 137 678 171
rect 626 99 678 137
rect 626 65 635 99
rect 669 65 678 99
rect 626 53 678 65
rect 712 387 764 399
rect 712 361 721 387
rect 755 361 764 387
rect 712 281 721 309
rect 755 281 764 309
rect 712 243 764 281
rect 712 209 721 243
rect 755 209 764 243
rect 712 171 764 209
rect 712 137 721 171
rect 755 137 764 171
rect 712 99 764 137
rect 712 65 721 99
rect 755 65 764 99
rect 712 53 764 65
rect 798 387 850 1365
rect 798 361 807 387
rect 841 361 850 387
rect 798 281 807 309
rect 841 281 850 309
rect 798 243 850 281
rect 798 209 807 243
rect 841 209 850 243
rect 798 171 850 209
rect 798 137 807 171
rect 841 137 850 171
rect 798 99 850 137
rect 798 65 807 99
rect 841 65 850 99
rect 798 53 850 65
<< via1 >>
rect 110 7537 162 7543
rect 110 7503 119 7537
rect 119 7503 153 7537
rect 153 7503 162 7537
rect 110 7491 162 7503
rect 196 7537 248 7543
rect 196 7503 205 7537
rect 205 7503 239 7537
rect 239 7503 248 7537
rect 196 7491 248 7503
rect 282 7537 334 7543
rect 282 7503 291 7537
rect 291 7503 325 7537
rect 325 7503 334 7537
rect 282 7491 334 7503
rect 196 6379 248 6409
rect 196 6357 205 6379
rect 205 6357 239 6379
rect 239 6357 248 6379
rect 368 7537 420 7543
rect 368 7503 377 7537
rect 377 7503 411 7537
rect 411 7503 420 7537
rect 368 7491 420 7503
rect 454 7537 506 7543
rect 454 7503 463 7537
rect 463 7503 497 7537
rect 497 7503 506 7537
rect 454 7491 506 7503
rect 540 7537 592 7543
rect 540 7503 549 7537
rect 549 7503 583 7537
rect 583 7503 592 7537
rect 540 7491 592 7503
rect 626 7537 678 7543
rect 626 7503 635 7537
rect 635 7503 669 7537
rect 669 7503 678 7537
rect 626 7491 678 7503
rect 398 6934 450 6986
rect 510 6934 562 6986
rect 196 5979 248 6031
rect 196 5246 248 5275
rect 196 5223 205 5246
rect 205 5223 239 5246
rect 239 5223 248 5246
rect 196 4845 248 4897
rect 196 4089 248 4141
rect 110 3099 162 3133
rect 110 3081 119 3099
rect 119 3081 153 3099
rect 153 3081 162 3099
rect 196 3315 248 3322
rect 196 3281 205 3315
rect 205 3281 239 3315
rect 239 3281 248 3315
rect 196 3270 248 3281
rect 282 3099 334 3133
rect 282 3081 291 3099
rect 291 3081 325 3099
rect 325 3081 334 3099
rect 196 2938 248 2944
rect 196 2904 205 2938
rect 205 2904 239 2938
rect 239 2904 248 2938
rect 196 2892 248 2904
rect 196 2514 248 2566
rect 196 1911 205 1936
rect 205 1911 239 1936
rect 239 1911 248 1936
rect 196 1884 248 1911
rect 398 2514 450 2566
rect 712 7537 764 7543
rect 712 7503 721 7537
rect 721 7503 755 7537
rect 755 7503 764 7537
rect 712 7491 764 7503
rect 798 7537 850 7543
rect 798 7503 807 7537
rect 807 7503 841 7537
rect 841 7503 850 7537
rect 798 7491 850 7503
rect 712 6379 764 6409
rect 712 6357 721 6379
rect 721 6357 755 6379
rect 755 6357 764 6379
rect 712 5979 764 6031
rect 712 5246 764 5275
rect 712 5223 721 5246
rect 721 5223 755 5246
rect 755 5223 764 5246
rect 712 4845 764 4897
rect 712 4089 764 4141
rect 712 3677 764 3700
rect 712 3648 721 3677
rect 721 3648 755 3677
rect 755 3648 764 3677
rect 510 2325 562 2377
rect 626 3099 678 3133
rect 626 3081 635 3099
rect 635 3081 669 3099
rect 669 3081 678 3099
rect 798 3099 850 3133
rect 798 3081 807 3099
rect 807 3081 841 3099
rect 841 3081 850 3099
rect 712 2938 764 2944
rect 712 2904 721 2938
rect 721 2904 755 2938
rect 755 2904 764 2938
rect 712 2892 764 2904
rect 712 2325 764 2377
rect 712 1911 721 1936
rect 721 1911 755 1936
rect 755 1911 764 1936
rect 712 1884 764 1911
rect 196 1238 248 1243
rect 196 1204 205 1238
rect 205 1204 239 1238
rect 239 1204 248 1238
rect 196 1191 248 1204
rect 110 353 119 361
rect 119 353 153 361
rect 153 353 162 361
rect 110 315 162 353
rect 110 309 119 315
rect 119 309 153 315
rect 153 309 162 315
rect 196 353 205 361
rect 205 353 239 361
rect 239 353 248 361
rect 196 315 248 353
rect 196 309 205 315
rect 205 309 239 315
rect 239 309 248 315
rect 282 353 291 361
rect 291 353 325 361
rect 325 353 334 361
rect 282 315 334 353
rect 282 309 291 315
rect 291 309 325 315
rect 325 309 334 315
rect 368 353 377 361
rect 377 353 411 361
rect 411 353 420 361
rect 368 315 420 353
rect 368 309 377 315
rect 377 309 411 315
rect 411 309 420 315
rect 454 353 463 361
rect 463 353 497 361
rect 497 353 506 361
rect 454 315 506 353
rect 454 309 463 315
rect 463 309 497 315
rect 497 309 506 315
rect 540 353 549 361
rect 549 353 583 361
rect 583 353 592 361
rect 540 315 592 353
rect 540 309 549 315
rect 549 309 583 315
rect 583 309 592 315
rect 712 1238 764 1243
rect 712 1204 721 1238
rect 721 1204 755 1238
rect 755 1204 764 1238
rect 712 1191 764 1204
rect 626 353 635 361
rect 635 353 669 361
rect 669 353 678 361
rect 626 315 678 353
rect 626 309 635 315
rect 635 309 669 315
rect 669 309 678 315
rect 712 353 721 361
rect 721 353 755 361
rect 755 353 764 361
rect 712 315 764 353
rect 712 309 721 315
rect 721 309 755 315
rect 755 309 764 315
rect 798 353 807 361
rect 807 353 841 361
rect 841 353 850 361
rect 798 315 850 353
rect 798 309 807 315
rect 807 309 841 315
rect 841 309 850 315
<< metal2 >>
rect 104 7543 856 7545
rect 104 7491 110 7543
rect 162 7491 196 7543
rect 248 7491 282 7543
rect 334 7491 368 7543
rect 420 7491 454 7543
rect 506 7491 540 7543
rect 592 7491 626 7543
rect 678 7491 712 7543
rect 764 7491 798 7543
rect 850 7491 856 7543
rect 104 7489 856 7491
rect 368 6988 456 6997
rect 368 6932 377 6988
rect 433 6986 456 6988
rect 450 6934 456 6986
rect 433 6932 456 6934
rect 368 6923 456 6932
rect 504 6988 592 6997
rect 504 6986 527 6988
rect 504 6934 510 6986
rect 504 6932 527 6934
rect 583 6932 592 6988
rect 504 6923 592 6932
rect 190 6409 366 6411
rect 190 6357 196 6409
rect 248 6357 366 6409
rect 190 6355 366 6357
rect 422 6355 431 6411
rect 529 6355 538 6411
rect 594 6409 770 6411
rect 594 6357 712 6409
rect 764 6357 770 6409
rect 594 6355 770 6357
rect 56 5977 65 6033
rect 121 6031 254 6033
rect 121 5979 196 6031
rect 248 5979 254 6031
rect 121 5977 254 5979
rect 706 6031 839 6033
rect 706 5979 712 6031
rect 764 5979 839 6031
rect 706 5977 839 5979
rect 895 5977 904 6033
rect 56 5221 65 5277
rect 121 5275 254 5277
rect 121 5223 196 5275
rect 248 5223 254 5275
rect 121 5221 254 5223
rect 706 5275 839 5277
rect 706 5223 712 5275
rect 764 5223 839 5275
rect 706 5221 839 5223
rect 895 5221 904 5277
rect 185 4843 194 4899
rect 250 4843 259 4899
rect 701 4843 710 4899
rect 766 4843 775 4899
rect 185 4087 194 4143
rect 250 4087 259 4143
rect 701 4087 710 4143
rect 766 4087 775 4143
rect 185 3646 194 3702
rect 250 3700 770 3702
rect 250 3648 712 3700
rect 764 3648 770 3700
rect 250 3646 770 3648
rect 190 3322 710 3324
rect 190 3270 196 3322
rect 248 3270 710 3322
rect 190 3268 710 3270
rect 766 3268 775 3324
rect 104 3133 366 3135
rect 104 3081 110 3133
rect 162 3081 282 3133
rect 334 3081 366 3133
rect 104 3079 366 3081
rect 422 3079 431 3135
rect 529 3079 538 3135
rect 594 3133 856 3135
rect 594 3081 626 3133
rect 678 3081 798 3133
rect 850 3081 856 3133
rect 594 3079 856 3081
rect 185 2890 194 2946
rect 250 2890 259 2946
rect 701 2890 710 2946
rect 766 2890 775 2946
rect 190 2566 770 2568
rect 190 2514 196 2566
rect 248 2514 398 2566
rect 450 2514 770 2566
rect 190 2512 770 2514
rect 190 2377 770 2379
rect 190 2325 510 2377
rect 562 2325 712 2377
rect 764 2325 770 2377
rect 190 2323 770 2325
rect 190 1936 770 1938
rect 190 1884 196 1936
rect 248 1884 712 1936
rect 764 1884 770 1936
rect 190 1882 770 1884
rect 56 1189 65 1245
rect 121 1243 839 1245
rect 121 1191 196 1243
rect 248 1191 712 1243
rect 764 1191 839 1243
rect 121 1189 839 1191
rect 895 1189 904 1245
rect 104 361 856 363
rect 104 309 110 361
rect 162 309 196 361
rect 248 309 282 361
rect 334 309 368 361
rect 420 309 454 361
rect 506 309 540 361
rect 592 309 626 361
rect 678 309 712 361
rect 764 309 798 361
rect 850 309 856 361
rect 104 307 856 309
<< via2 >>
rect 377 6986 433 6988
rect 377 6934 398 6986
rect 398 6934 433 6986
rect 377 6932 433 6934
rect 527 6986 583 6988
rect 527 6934 562 6986
rect 562 6934 583 6986
rect 527 6932 583 6934
rect 366 6355 422 6411
rect 538 6355 594 6411
rect 65 5977 121 6033
rect 839 5977 895 6033
rect 65 5221 121 5277
rect 839 5221 895 5277
rect 194 4897 250 4899
rect 194 4845 196 4897
rect 196 4845 248 4897
rect 248 4845 250 4897
rect 194 4843 250 4845
rect 710 4897 766 4899
rect 710 4845 712 4897
rect 712 4845 764 4897
rect 764 4845 766 4897
rect 710 4843 766 4845
rect 194 4141 250 4143
rect 194 4089 196 4141
rect 196 4089 248 4141
rect 248 4089 250 4141
rect 194 4087 250 4089
rect 710 4141 766 4143
rect 710 4089 712 4141
rect 712 4089 764 4141
rect 764 4089 766 4141
rect 710 4087 766 4089
rect 194 3646 250 3702
rect 710 3268 766 3324
rect 366 3079 422 3135
rect 538 3079 594 3135
rect 194 2944 250 2946
rect 194 2892 196 2944
rect 196 2892 248 2944
rect 248 2892 250 2944
rect 194 2890 250 2892
rect 710 2944 766 2946
rect 710 2892 712 2944
rect 712 2892 764 2944
rect 764 2892 766 2944
rect 710 2890 766 2892
rect 65 1189 121 1245
rect 839 1189 895 1245
<< metal3 >>
rect 368 6988 442 7737
rect 368 6932 377 6988
rect 433 6932 442 6988
rect 368 6925 442 6932
rect 518 6988 592 7737
rect 518 6932 527 6988
rect 583 6932 592 6988
rect 518 6925 592 6932
rect 361 6411 427 6420
rect 361 6355 366 6411
rect 422 6355 427 6411
rect 60 6033 126 6042
rect 60 5977 65 6033
rect 121 5977 126 6033
rect 60 5277 126 5977
rect 60 5221 65 5277
rect 121 5221 126 5277
rect 60 1245 126 5221
rect 189 4899 255 4908
rect 189 4843 194 4899
rect 250 4843 255 4899
rect 189 4143 255 4843
rect 189 4087 194 4143
rect 250 4087 255 4143
rect 189 3702 255 4087
rect 189 3646 194 3702
rect 250 3646 255 3702
rect 189 2946 255 3646
rect 361 3135 427 6355
rect 361 3079 366 3135
rect 422 3079 427 3135
rect 361 3070 427 3079
rect 533 6411 599 6420
rect 533 6355 538 6411
rect 594 6355 599 6411
rect 533 3135 599 6355
rect 834 6033 900 6042
rect 834 5977 839 6033
rect 895 5977 900 6033
rect 834 5277 900 5977
rect 834 5221 839 5277
rect 895 5221 900 5277
rect 533 3079 538 3135
rect 594 3079 599 3135
rect 533 3070 599 3079
rect 705 4899 771 4908
rect 705 4843 710 4899
rect 766 4843 771 4899
rect 705 4143 771 4843
rect 705 4087 710 4143
rect 766 4087 771 4143
rect 705 3324 771 4087
rect 705 3268 710 3324
rect 766 3268 771 3324
rect 189 2890 194 2946
rect 250 2890 255 2946
rect 189 2881 255 2890
rect 705 2946 771 3268
rect 705 2890 710 2946
rect 766 2890 771 2946
rect 705 2881 771 2890
rect 60 1189 65 1245
rect 121 1189 126 1245
rect 60 1180 126 1189
rect 834 1245 900 5221
rect 834 1189 839 1245
rect 895 1189 900 1245
rect 834 1180 900 1189
<< labels >>
flabel metal2 104 307 856 363 0 FreeSans 560 0 0 0 sa_senseamp_0/VSS
flabel metal2 104 7489 856 7545 0 FreeSans 560 0 0 0 sa_senseamp_0/VDD
flabel metal2 190 1189 770 1245 0 FreeSans 560 0 0 0 sa_senseamp_0/clk
flabel metal2 190 2323 770 2379 0 FreeSans 560 0 0 0 sa_senseamp_0/inn
flabel metal2 190 2512 770 2568 0 FreeSans 560 0 0 0 sa_senseamp_0/inp
flabel metal3 705 2881 771 4908 0 FreeSans 660 90 0 0 sa_senseamp_0/outn
flabel metal3 189 2881 255 4908 0 FreeSans 660 90 0 0 sa_senseamp_0/outp
flabel metal3 361 3070 427 6420 0 FreeSans 660 90 0 0 sa_senseamp_0/midn
flabel metal3 533 3070 599 6420 0 FreeSans 660 90 0 0 sa_senseamp_0/midp
<< end >>
