.SUBCKT dbdr_nand
+ a b y vdd gnd

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dbdr_inv 
+ din din_b vdd gnd

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.subckt dbdr_delay_cell clk_in clk_out en din dout vdd vss
Xinv clk_in int vdd vss dbdr_inv
Xnand_clk int din clk_out vdd vss dbdr_nand
Xnand_out int en dout vdd vss dbdr_nand
.ends
