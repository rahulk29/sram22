.subckt dbdr_delay_unit_3 clk_in clk_out sae_in sae_out clk_rev vdd vss
X0 clk_in clk_out sae_in vdd nn vdd vss dbdr_delay_cell
X1 clk_rev int12 vdd nn noconn0 vdd vss dbdr_delay_cell
X2 int12 sae_out vdd vdd noconn1 vdd vss dbdr_delay_cell
.ends

.subckt timing_multiplier_3 clk sae_in sae_out vdd vss
X0 clk f0 sae_in sae_out clk_rev_0 vdd vss dbdr_delay_unit_3
X1 f0 f1 sae_in clk_rev_0 clk_rev_1 vdd vss dbdr_delay_unit_3
X2 f1 f2 sae_in clk_rev_1 clk_rev_2 vdd vss dbdr_delay_unit_3
X3 f2 f3 sae_in clk_rev_2 clk_rev_3 vdd vss dbdr_delay_unit_3
X4 f3 f4 sae_in clk_rev_3 clk_rev_4 vdd vss dbdr_delay_unit_3
X5 f4 f5 sae_in clk_rev_4 clk_rev_5 vdd vss dbdr_delay_unit_3
X6 f5 f6 sae_in clk_rev_5 clk_rev_6 vdd vss dbdr_delay_unit_3
X7 f6 f7 sae_in clk_rev_6 clk_rev_7 vdd vss dbdr_delay_unit_3
X8 f7 f8 sae_in clk_rev_7 clk_rev_8 vdd vss dbdr_delay_unit_3
X9 f8 f9 sae_in clk_rev_8 clk_rev_9 vdd vss dbdr_delay_unit_3
X10 f9 f10 sae_in clk_rev_9 clk_rev_10 vdd vss dbdr_delay_unit_3
X11 f10 f11 sae_in clk_rev_10 clk_rev_11 vdd vss dbdr_delay_unit_3
X12 f11 f12 sae_in clk_rev_11 clk_rev_12 vdd vss dbdr_delay_unit_3
X13 f12 f13 sae_in clk_rev_12 clk_rev_13 vdd vss dbdr_delay_unit_3
X14 f13 f14 sae_in clk_rev_13 clk_rev_14 vdd vss dbdr_delay_unit_3
X15 f14 f15 sae_in clk_rev_14 clk_rev_15 vdd vss dbdr_delay_unit_3
X16 f15 f16 sae_in clk_rev_15 clk_rev_16 vdd vss dbdr_delay_unit_3
X17 f16 f17 sae_in clk_rev_16 clk_rev_17 vdd vss dbdr_delay_unit_3
X18 f17 f18 sae_in clk_rev_17 clk_rev_18 vdd vss dbdr_delay_unit_3
X19 f18 f19 sae_in clk_rev_18 clk_rev_19 vdd vss dbdr_delay_unit_3
X20 f19 f20 sae_in clk_rev_19 vss vdd vss dbdr_delay_unit_3
.ends
