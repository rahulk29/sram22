* empty netlist
