* Voltage divider

V1 in 0 dc 1
R1 in out 1k
R2 out 0 1k

.end
