magic
tech sky130A
magscale 1 2
timestamp 1644438400
<< nwell >>
rect 168 0 548 316
<< nmos >>
rect -100 186 100 216
rect -100 100 100 130
<< pmos >>
rect 204 186 512 216
rect 204 100 512 130
<< ndiff >>
rect -100 261 100 269
rect -100 227 -51 261
rect -17 227 17 261
rect 51 227 100 261
rect -100 216 100 227
rect -100 175 100 186
rect -100 141 -51 175
rect -17 141 17 175
rect 51 141 100 175
rect -100 130 100 141
rect -100 89 100 100
rect -100 55 -51 89
rect -17 55 17 89
rect 51 55 100 89
rect -100 47 100 55
<< pdiff >>
rect 204 261 512 269
rect 204 227 239 261
rect 273 227 307 261
rect 341 227 375 261
rect 409 227 443 261
rect 477 227 512 261
rect 204 216 512 227
rect 204 175 512 186
rect 204 141 239 175
rect 273 141 307 175
rect 341 141 375 175
rect 409 141 443 175
rect 477 141 512 175
rect 204 130 512 141
rect 204 89 512 100
rect 204 55 239 89
rect 273 55 307 89
rect 341 55 375 89
rect 409 55 443 89
rect 477 55 512 89
rect 204 47 512 55
<< ndiffc >>
rect -51 227 -17 261
rect 17 227 51 261
rect -51 141 -17 175
rect 17 141 51 175
rect -51 55 -17 89
rect 17 55 51 89
<< pdiffc >>
rect 239 227 273 261
rect 307 227 341 261
rect 375 227 409 261
rect 443 227 477 261
rect 239 141 273 175
rect 307 141 341 175
rect 375 141 409 175
rect 443 141 477 175
rect 239 55 273 89
rect 307 55 341 89
rect 375 55 409 89
rect 443 55 477 89
<< poly >>
rect -192 230 -126 240
rect -192 196 -176 230
rect -142 216 -126 230
rect -142 196 -100 216
rect -192 186 -100 196
rect 100 186 204 216
rect 512 186 538 216
rect -192 120 -100 130
rect -192 86 -176 120
rect -142 100 -100 120
rect 100 100 204 130
rect 512 100 538 130
rect -142 86 -126 100
rect -192 76 -126 86
<< polycont >>
rect -176 196 -142 230
rect -176 86 -142 120
<< locali >>
rect -176 230 -142 246
rect -100 227 -51 261
rect 51 227 100 261
rect 204 227 239 261
rect 273 227 307 261
rect 409 227 443 261
rect 477 227 512 261
rect -176 120 -142 196
rect -100 141 -51 175
rect -17 141 17 175
rect 51 141 239 175
rect 273 141 307 175
rect 341 141 375 175
rect 409 141 443 175
rect 477 141 512 175
rect -176 70 -142 86
rect -100 55 -51 89
rect 51 55 100 89
rect 204 55 239 89
rect 273 55 307 89
rect 409 55 443 89
rect 477 55 512 89
<< viali >>
rect -17 227 17 261
rect 341 227 375 261
rect -17 55 17 89
rect 341 55 375 89
<< metal1 >>
rect -192 299 548 316
rect -29 261 29 267
rect -29 227 -17 261
rect 17 227 29 261
rect -29 89 29 227
rect -29 55 -17 89
rect 17 55 29 89
rect -29 17 29 55
rect 329 261 387 299
rect 329 227 341 261
rect 375 227 387 261
rect 329 89 387 227
rect 329 55 341 89
rect 375 55 387 89
rect 329 49 387 55
rect -192 0 548 17
<< labels >>
rlabel nwell 168 0 548 316 3 VPB
port 3 e
rlabel locali -100 141 512 175 3 Y
port 5 e
rlabel locali -176 70 -142 246 7 A
port 0 w
rlabel metal1 -192 299 548 316 7 VPWR
port 4 w
rlabel metal1 -192 0 548 17 7 VGND
port 1 w
<< end >>
