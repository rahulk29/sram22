magic
tech sky130A
magscale 1 2
timestamp 1645319861
<< checkpaint >>
rect -1000 1487 1552 1508
rect -1294 -1147 1552 1487
rect -1294 -1169 1260 -1147
<< dnwell >>
rect 0 0 260 316
<< pwell >>
rect 57 200 203 278
rect 0 116 260 200
rect 57 96 203 116
<< ndiff >>
rect 14 142 27 174
rect 233 142 246 174
<< ndiffc >>
rect 0 142 14 174
rect 246 142 260 174
<< psubdiff >>
rect 83 245 177 252
rect 83 211 113 245
rect 147 211 177 245
rect 83 177 177 211
rect 83 143 113 177
rect 147 143 177 177
rect 83 122 177 143
<< psubdiffcont >>
rect 113 211 147 245
rect 113 143 147 177
<< poly >>
rect 0 262 260 292
rect 40 90 73 262
rect 187 90 220 262
rect 40 74 220 90
rect 40 54 56 74
rect 0 40 56 54
rect 90 40 170 74
rect 204 54 220 74
rect 204 40 260 54
rect 0 24 260 40
<< polycont >>
rect 56 40 90 74
rect 170 40 204 74
<< corelocali >>
rect 44 211 113 245
rect 147 227 216 245
rect 147 211 165 227
rect 44 193 165 211
rect 199 193 216 227
rect 0 175 14 191
rect 44 177 216 193
rect 44 143 113 177
rect 147 155 216 177
rect 246 175 260 191
rect 147 143 165 155
rect 0 125 14 141
rect 44 121 165 143
rect 199 121 216 155
rect 246 125 260 141
rect 44 107 216 121
rect 40 40 56 74
rect 90 66 170 74
rect 90 40 113 66
rect 147 40 170 66
rect 204 40 220 74
<< viali >>
rect 165 193 199 227
rect 0 174 17 175
rect 0 142 14 174
rect 14 142 17 174
rect 0 141 17 142
rect 165 121 199 155
rect 243 174 260 175
rect 243 142 246 174
rect 246 142 260 174
rect 243 141 260 142
rect 113 32 147 66
<< metal1 >>
rect 0 263 14 316
rect 0 178 26 263
rect 25 128 26 178
rect 0 126 26 128
rect 0 121 21 126
tri 21 121 26 126 nw
rect 0 0 14 121
rect 54 116 102 316
tri 42 102 54 114 se
rect 54 102 76 116
rect 42 0 76 102
tri 76 90 102 116 nw
rect 158 227 206 316
rect 246 263 260 316
rect 158 193 165 227
rect 199 193 206 227
rect 158 155 206 193
rect 158 121 165 155
rect 199 121 206 155
rect 234 178 260 263
rect 234 128 235 178
rect 234 126 260 128
tri 234 121 239 126 ne
rect 239 121 260 126
rect 158 116 206 121
tri 158 90 184 116 ne
rect 184 102 206 116
tri 206 102 218 114 sw
tri 104 75 111 82 se
rect 111 75 149 82
tri 149 75 156 82 sw
rect 104 74 156 75
rect 104 24 105 74
rect 155 24 156 74
rect 104 21 156 24
tri 104 14 111 21 ne
rect 111 14 149 21
tri 149 14 156 21 nw
rect 184 0 218 102
rect 246 0 260 121
<< via1 >>
rect 0 175 25 178
rect 0 141 17 175
rect 17 141 25 175
rect 0 128 25 141
rect 235 175 260 178
rect 235 141 243 175
rect 243 141 260 175
rect 235 128 260 141
rect 105 66 155 74
rect 105 32 113 66
rect 113 32 147 66
rect 147 32 155 66
rect 105 24 155 32
<< metal2 >>
rect 0 213 260 257
rect 0 178 260 179
rect 25 128 235 178
rect 0 127 260 128
rect 0 74 260 93
rect 0 59 105 74
rect 98 24 105 59
rect 155 59 260 74
rect 155 24 162 59
<< labels >>
rlabel metal1 s 0 0 14 15 4 VGND
rlabel metal1 s 246 0 260 15 4 VGND
<< end >>
