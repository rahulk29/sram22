************************************************************************
* auCdl Netlist:
* 
* Library Name:  AAA_Comp_SA_layers
* Top Cell Name: AAA_Comp_SA_sense
* View Name:     schematic
* Netlisted on:  Nov  1 17:24:53 2022
************************************************************************
*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
* .PARAM
************************************************************************
* Library Name: BAG_prim
* Cell Name:    nmos4_standard_pcell_0
* View Name:    schematic
************************************************************************
.SUBCKT nmos4_standard_pcell_0 B D G S
*.PININFO B:B D:B G:B S:B
XN0 D G S B sky130_fd_pr__nfet_01v8 m=4 w=1.68 l=0.15 mult=1 sa=0.0 sb=0.0 sd=0.0 
+ topography=normal area=0.063 perim=1.14
.ENDS
************************************************************************
* Library Name: BAG_prim
* Cell Name:    nmos4_standard_pcell_1
* View Name:    schematic
************************************************************************
.SUBCKT nmos4_standard_pcell_1 B D G S
*.PININFO B:B D:B G:B S:B
XN0 D G S B sky130_fd_pr__nfet_01v8 m=2 w=1.68 l=0.15 mult=1 sa=0.0 sb=0.0 sd=0.0 
+ topography=normal area=0.063 perim=1.14
.ENDS
************************************************************************
* Library Name: BAG_prim
* Cell Name:    pmos4_standard_pcell_2
* View Name:    schematic
************************************************************************
.SUBCKT pmos4_standard_pcell_2 B D G S
*.PININFO B:B D:B G:B S:B
XN0 D G S B sky130_fd_pr__pfet_01v8 m=2 w=1.00 l=0.15 mult=1 sa=0.0 sb=0.0 sd=0.0 
+ topography=normal area=0.063 perim=1.14
.ENDS
************************************************************************
* Library Name: BAG_prim
* Cell Name:    pmos4_standard_pcell_3
* View Name:    schematic
************************************************************************
.SUBCKT pmos4_standard_pcell_3 B D G S
*.PININFO B:B D:B G:B S:B
XN0 D G S B sky130_fd_pr__pfet_01v8 m=2 w=2.00 l=0.15 mult=1 sa=0.0 sb=0.0 sd=0.0 
+ topography=normal area=0.063 perim=1.14
.ENDS
************************************************************************
* Library Name: AAA_Comp_SA_layers
* Cell Name:    AAA_Comp_SA_sense
* View Name:    schematic
************************************************************************
.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS
*.PININFO clk:I inn:I inp:I midn:O midp:O outn:O outp:O VDD:B VSS:B
XXTAIL VSS tail clk VSS nmos4_standard_pcell_0
XXNFBP VSS outp outn midp nmos4_standard_pcell_1
XXNFBN VSS outn outp midn nmos4_standard_pcell_1
XXINP VSS midn inp tail nmos4_standard_pcell_1
XXINN VSS midp inn tail nmos4_standard_pcell_1
XXSWOP VDD outp clk VDD pmos4_standard_pcell_2
XXSWON VDD outn clk VDD pmos4_standard_pcell_2
XXSWMP VDD midp clk VDD pmos4_standard_pcell_2
XXSWMN VDD midn clk VDD pmos4_standard_pcell_2
XXPFBP VDD outp outn VDD pmos4_standard_pcell_3
XXPFBN VDD outn outp VDD pmos4_standard_pcell_3
.ENDS
