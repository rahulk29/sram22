magic
tech sky130A
timestamp 1643225352
<< nwell >>
rect 460 0 605 105
<< pwell >>
rect 469 -112 554 -27
rect 504 -117 519 -112
<< nmos >>
rect 504 -102 519 -37
<< pmos >>
rect 505 20 520 85
rect 545 20 560 85
<< ndiff >>
rect 479 -102 504 -37
rect 519 -102 544 -37
<< pdiff >>
rect 480 20 505 85
rect 520 20 545 85
rect 560 20 585 85
<< poly >>
rect 505 85 520 105
rect 545 85 560 105
rect 505 0 520 20
rect 545 0 560 20
rect 504 -37 519 -22
rect 504 -117 519 -102
<< metal2 >>
rect 670 -91 790 67
<< properties >>
string FIXED_BBOX 0 0 138 272
string path 0.000 0.000 2.760 0.000 
<< end >>
