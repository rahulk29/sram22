magic
tech sky130A
magscale 1 2
timestamp 1644441317
<< checkpaint >>
rect -1260 -1260 2000 1587
<< locali >>
rect 0 227 50 261
rect 0 55 50 89
use inv_pm_sh_2  inv_pm_sh_2_0 ~/acads/sky130/sram22/tech/sky130/magic
timestamp 1644438400
transform 1 0 192 0 1 0
box -192 0 548 316
use wl_route  wl_route_0 ~/acads/sky130/sram22/tech/sky130/magic
timestamp 1644435965
transform 1 0 753 0 1 282
box -151 -232 -13 -101
<< end >>
