magic
tech sky130A
timestamp 1644438400
<< nwell >>
rect 84 0 274 158
<< nmos >>
rect -50 93 50 108
rect -50 50 50 65
<< pmos >>
rect 102 93 256 108
rect 102 50 256 65
<< ndiff >>
rect -50 130 50 134
rect -50 113 -25 130
rect -8 113 8 130
rect 25 113 50 130
rect -50 108 50 113
rect -50 87 50 93
rect -50 70 -25 87
rect -8 70 8 87
rect 25 70 50 87
rect -50 65 50 70
rect -50 44 50 50
rect -50 27 -25 44
rect -8 27 8 44
rect 25 27 50 44
rect -50 23 50 27
<< pdiff >>
rect 102 130 256 134
rect 102 113 119 130
rect 136 113 153 130
rect 170 113 187 130
rect 204 113 221 130
rect 238 113 256 130
rect 102 108 256 113
rect 102 87 256 93
rect 102 70 119 87
rect 136 70 153 87
rect 170 70 187 87
rect 204 70 221 87
rect 238 70 256 87
rect 102 65 256 70
rect 102 44 256 50
rect 102 27 119 44
rect 136 27 153 44
rect 170 27 187 44
rect 204 27 221 44
rect 238 27 256 44
rect 102 23 256 27
<< ndiffc >>
rect -25 113 -8 130
rect 8 113 25 130
rect -25 70 -8 87
rect 8 70 25 87
rect -25 27 -8 44
rect 8 27 25 44
<< pdiffc >>
rect 119 113 136 130
rect 153 113 170 130
rect 187 113 204 130
rect 221 113 238 130
rect 119 70 136 87
rect 153 70 170 87
rect 187 70 204 87
rect 221 70 238 87
rect 119 27 136 44
rect 153 27 170 44
rect 187 27 204 44
rect 221 27 238 44
<< poly >>
rect -96 115 -63 120
rect -96 98 -88 115
rect -71 108 -63 115
rect -71 98 -50 108
rect -96 93 -50 98
rect 50 93 102 108
rect 256 93 269 108
rect -96 60 -50 65
rect -96 43 -88 60
rect -71 50 -50 60
rect 50 50 102 65
rect 256 50 269 65
rect -71 43 -63 50
rect -96 38 -63 43
<< polycont >>
rect -88 98 -71 115
rect -88 43 -71 60
<< locali >>
rect -88 115 -71 123
rect -50 113 -25 130
rect 25 113 50 130
rect 102 113 119 130
rect 136 113 153 130
rect 204 113 221 130
rect 238 113 256 130
rect -88 60 -71 98
rect -50 70 -25 87
rect -8 70 8 87
rect 25 70 119 87
rect 136 70 153 87
rect 170 70 187 87
rect 204 70 221 87
rect 238 70 256 87
rect -88 35 -71 43
rect -50 27 -25 44
rect 25 27 50 44
rect 102 27 119 44
rect 136 27 153 44
rect 204 27 221 44
rect 238 27 256 44
<< viali >>
rect -8 113 8 130
rect 170 113 187 130
rect -8 27 8 44
rect 170 27 187 44
<< metal1 >>
rect -96 149 274 158
rect -14 130 14 133
rect -14 113 -8 130
rect 8 113 14 130
rect -14 44 14 113
rect -14 27 -8 44
rect 8 27 14 44
rect -14 8 14 27
rect 164 130 193 149
rect 164 113 170 130
rect 187 113 193 130
rect 164 44 193 113
rect 164 27 170 44
rect 187 27 193 44
rect 164 24 193 27
rect -96 0 274 8
<< labels >>
rlabel nwell 84 0 274 158 3 VPB
port 3 e
rlabel locali -50 70 256 87 3 Y
port 5 e
rlabel locali -88 35 -71 123 7 A
port 0 w
rlabel metal1 -96 149 274 158 7 VPWR
port 4 w
rlabel metal1 -96 0 274 8 7 VGND
port 1 w
<< end >>
