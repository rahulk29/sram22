* Sramgen control circuit

.subckt control_logic_inv0 din din_b vdd vss
Xp din_b din vdd vdd sky130_fd_pr__pfet_01v8 w='1' l='0.15'
Xn din_b din vss vss sky130_fd_pr__nfet_01v8 w='0.6' l='0.15'
.ends

.subckt control_logic_delay_chain din din_b dout vdd vss
Xinv0 din din_b vdd vss control_logic_inv0
Xinv1 din_b tmp1 vdd vss control_logic_inv0
Xinv2 tmp1 tmp2 vdd vss control_logic_inv0
Xinv3 tmp2 tmp3 vdd vss control_logic_inv0
Xinv4 tmp3 tmp4 vdd vss control_logic_inv0
Xinv5 tmp4 tmp5 vdd vss control_logic_inv0
Xinv6 tmp5 tmp6 vdd vss control_logic_inv0
Xinv7 tmp6 tmp7 vdd vss control_logic_inv0
Xinv8 tmp7 tmp8 vdd vss control_logic_inv0
Xinv9 tmp8 tmp9 vdd vss control_logic_inv0
Xinv10 tmp9 tmp10 vdd vss control_logic_inv0
Xinv11 tmp10 tmp11 vdd vss control_logic_inv0
Xinv12 tmp11 tmp12 vdd vss control_logic_inv0
Xinv13 tmp12 tmp13 vdd vss control_logic_inv0
Xinv14 tmp13 tmp14 vdd vss control_logic_inv0
Xinv15 tmp14 dout vdd vss control_logic_inv0
.ends

.subckt control_logic_nand0 a b y vdd vss
Xp1 y a vdd vdd sky130_fd_pr__pfet_01v8 w='2' l='0.15'
Xp2 y b vdd vdd sky130_fd_pr__pfet_01v8 w='2' l='0.15'
Xn1 y a int vss sky130_fd_pr__nfet_01v8 w='1' l='0.15'
Xn2 int b vss vss sky130_fd_pr__nfet_01v8 w='1' l='0.15'
.ends

.subckt control_logic_and0 a b y vdd vss
Xnand a b y_bar vdd vss control_logic_nand0
Xinv y_bar y vdd vss control_logic_inv0
.ends

.subckt control_logic_nor a b y vdd vss
* Y = !(A || B)
Xn1 y a vss vss sky130_fd_pr__nfet_01v8 w='1' l='0.15'
Xn2 y b vss vss sky130_fd_pr__nfet_01v8 w='1' l='0.15'
Xp1 int a vdd vdd sky130_fd_pr__pfet_01v8 w='3' l='0.15'
Xp2 y b int vdd sky130_fd_pr__pfet_01v8 w='3' l='0.15'
.ends

.subckt control_logic_sr_latch set reset q q_b vdd vss
Xnor1 set q q_b vdd vss control_logic_nor
Xnor2 reset q_b q vdd vss control_logic_nor
.ends

.subckt sramgen_control clk cs we sae_i pc pc_b wl_en write_driver_en sense_en vdd vss
* INPUT: clk cs we sae_i
* OUTPUT: pc pc_b wl_en write_driver_en sense_en
* INOUT: vdd vss

* PC = CLK && CS
Xand0 clk cs pc vdd vss control_logic_and0

* PC_B = !PC
Xinv_pc pc pc_b vdd vss control_logic_inv0

* CLK_B = !CLK
Xinv_clk clk clk_b vdd vss control_logic_inv0

* CLK_B_GATED = CLK_B && CS
Xand1 clk_b cs clk_b_gated vdd vss control_logic_and0

* WRITE_DRIVER_EN = CLK_B_GATED && WE
Xand2 clk_b_gated we write_driver_en vdd vss control_logic_and0

* WL_EN = delay(CLK_B_GATED)
Xdelay_wl_en clk_b_gated clk_b_gated_b wl_en vdd vss control_logic_delay_chain

* SAE_O = delay WL_EN by 3 times T(sae_i) - T(wl_en)
Xtmc wl_en sae_i sae_o vdd vss timing_multiplier_3

* SENSE_EN = latched SAE_O
Xsae_latch sae_o clk sense_en sense_en_b vdd vss control_logic_sr_latch
.ends

