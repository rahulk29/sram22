* SRAM 16x16 simple READ testbench

.lib /Users/rahul/acads/research/sky130/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt

.include ../../lib/sram_sp_cell/sky130_fd_bd_sram__sram_sp_cell.spice
.include ../../lib/sramgen_control/sramgen_control.spice
.include ../../lib/sramgen_sp_sense_amp/sramgen_sp_sense_amp.spice

.include ../../build/ngspice/sram_16x16m2.spice

.param cload='20f'
.param vdd='1.8'
.param tr='10p'
.param tf='10p'

Xsram
+ vdd 0 clk
* din
+ vdd vdd vdd 0    vdd 0 vdd 0    0 vdd vdd vdd    vdd 0 0 vdd
* din_b
+ 0 0 0 vdd        0 vdd 0 vdd    vdd 0 0 0        0 vdd vdd 0
* dout
+ dout_3 dout_2 dout_1 dout_0
* we cs
+ 0 vdd
* addr
+ vdd 0 vdd 0 vdd 0
* addr_b
+ 0 vdd 0 vdd 0 vdd 
+ sramgen_sram_16x16m2

* 250 MHz clock
Vclk clk 0 dc 0 PULSE(0 {vdd} 10p {tr} {tf} 2n 4n 0)
Vdd vdd 0 {vdd}

Co1 dout_0 0 {cload}
Co2 dout_1 0 {cload}
Co3 dout_2 0 {cload}
Co4 dout_3 0 {cload}

.ic 
+ v(xsram.xbitcells.xbitcell_10_0.q)={vdd}
+ v(xsram.xbitcells.xbitcell_10_1.q)={vdd}
+ v(xsram.xbitcells.xbitcell_10_2.q)={vdd}
+ v(xsram.xbitcells.xbitcell_10_3.q)={vdd}
+ v(xsram.xbitcells.xbitcell_10_4.q)=0
+ v(xsram.xbitcells.xbitcell_10_5.q)=0
+ v(xsram.xbitcells.xbitcell_10_6.q)=0
+ v(xsram.xbitcells.xbitcell_10_7.q)=0
+ v(dout_3)=0
+ v(dout_2)=0
+ v(dout_1)=0
+ v(dout_0)=0

.control

tran 5p 12n 0u
wrdata read.dat
+ v(clk)
+ v(dout_3)
+ v(dout_2)
+ v(dout_1)
+ v(dout_0)
+ v(xsram.pc_b)
+ v(xsram.wl_en)
+ v(xsram.wr_drv_en)
+ v(xsram.xbitcells.xbitcell_10_0.q)
+ v(xsram.xbitcells.xbitcell_10_1.q)
+ v(xsram.xbitcells.xbitcell_10_2.q)
+ v(xsram.xbitcells.xbitcell_10_3.q)
+ v(xsram.xbitcells.xbitcell_10_4.q)
+ v(xsram.xbitcells.xbitcell_10_5.q)
+ v(xsram.xbitcells.xbitcell_10_6.q)
+ v(xsram.xbitcells.xbitcell_10_7.q)
unset askquit
quit 0
.endc

.end

