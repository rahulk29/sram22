* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell.ext - technology: sky130A

.subckt sram_sp_cell BL BR VDD VSS WL VNB VPB
X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass ad=0.04375 pd=0.92 as=0.0168 ps=0.52 w=0.14 l=0.15
X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch ad=0.156 pd=2.38 as=0.0808 ps=1.28 w=0.21 l=0.15
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass ad=0.0168 pd=0.52 as=0.0425 ps=0.92 w=0.14 l=0.15
X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass ad=0.064 pd=1.14 as=0p ps=0u w=0.14 l=0.15
X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=0.14 l=0.15
X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21 l=0.15
.ends

.subckt sky130_fd_bd_sram__sram_sp_colend BL1 VPWR VGND BL0 VNB VPB
.ends

