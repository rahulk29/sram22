* SRAM 4x4 read testbench

.lib /Users/rahul/acads/research/sky130/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice ff

.include ../../lib/sram_sp_cell/sky130_fd_bd_sram__sram_sp_cell.spice
.include ../../lib/sramgen_sp_sense_amp/sramgen_sp_sense_amp.spice
.include ../../lib/sramgen_control/sramgen_control_simple.spice
.include ../../lib/openram_dff/openram_dff.spice
.include ../../build/ngspice/sram_4x4m2.spice

.param vdd='1.8'
.param tr='100p'
.param tf='100p'


Xsram
* vdd vss clk 
+ vdd vss clk
* din_in_1 din_in_0
+ vss vss
* dout_1 dout_0
+ dout_1 dout_0
* we
+ we
* addr_in_2 addr_in_1 addr_in_0 
+ vdd vss vss
+ sramgen_sram_4x4m2

Vclk clk 0 dc 1.8 PULSE(0 {vdd} 10p {tr} {tf} 2n 4n 0)
Vss vss 0 dc 0
Vdd vdd 0 {vdd}
Vwe we 0 dc 1.8 PULSE({vdd} 0 0 {tr} {tf} 3n 100 0}

.ic
+ v(clk)=1.8
+ v(xsram.xbitcells.xbitcell_2_0.q)=1.8
+ v(xsram.xbitcells.xbitcell_2_0.qb)=0.0
+ v(xsram.xbitcells.xbitcell_2_2.q)=1.8
+ v(xsram.xbitcells.xbitcell_2_2.qb)=0.0
+ v(bl_0)=1.8
+ v(br_0)=1.8
+ v(bl_1)=1.8
+ v(br_1)=1.8
+ v(bl_2)=1.8
+ v(br_2)=1.8
+ v(bl_3)=1.8
+ v(br_3)=1.8

.control
tran 5p 18n 0n
wrdata read.dat
+ v(vdd)
+ v(vss)
+ v(clk)
+ v(dout_1)
+ v(dout_0)
+ v(xsram.wl_3)
+ v(xsram.wl_2)
+ v(xsram.wl_1)
+ v(xsram.wl_0)
+ v(xsram.bl_3)
+ v(xsram.bl_2)
+ v(xsram.bl_1)
+ v(xsram.bl_0)
+ v(xsram.br_3)
+ v(xsram.br_2)
+ v(xsram.br_1)
+ v(xsram.br_0)
+ v(xsram.bl_read_1)
+ v(xsram.br_read_1)
+ v(xsram.bl_read_0)
+ v(xsram.br_read_0)
+ v(xsram.bank_addr_0)
+ v(xsram.bank_addr_b_0)
+ v(xsram.sense_amp_en)
+ v(xsram.xsense_amp_array.data_b_0)
+ v(xsram.xbitcells.xbitcell_2_0.q)
+ v(xsram.xbitcells.xbitcell_2_0.qb)
.endc

.end

