* Sramgen control circuit

* Standard cells
* .subckt sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
.subckt control_logic_inv din din_b vdd vss
X0 vss din din_b vss sky130_fd_pr__nfet_01v8_lvt w=0.74 l=150000u
X1 din_b din vdd vdd sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 vdd din din_b vdd sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 din_b din vss vss sky130_fd_pr__nfet_01v8_lvt w=0.74 l=150000u
.ends

* .subckt sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X
.subckt control_logic_and2 A B X vdd vss
X0 a_31_74# B vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 X a_31_74# vss vss sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 X a_31_74# vdd vdd sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_118_74# B vss vss sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_31_74# A a_118_74# vss sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 vdd A a_31_74# vdd sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 vdd a_31_74# X vdd sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 vss a_31_74# X vss sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* .subckt sky130_fd_sc_hs__nor2_2 A B VGND VNB VPB VPWR Y
.subckt control_logic_nor2 A B Y VGND VNB VPB VPWR
X0 a_35_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_35_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y B a_35_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR A a_35_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* .subckt sky130_fd_sc_hs__or2_2 A B VGND VNB VPB VPWR X
.subckt control_logic_or2 A B X VPWR VGND
X0 VGND a_27_368# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_27_368# B a_114_368# VPWR sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 a_27_368# A VGND VGND sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND B a_27_368# VGND sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_114_368# A VPWR VPWR sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 X a_27_368# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 X a_27_368# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_27_368# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends

.SUBCKT control_logic_sr_latch 
+ s r q qb vdd vss 

xnor_set 
+ s q qb vss vss vdd vdd
+ control_logic_nor2 
* No parameters

xnor_reset 
+ r qb q vss vss vdd vdd
+ control_logic_nor2 
* No parameters

.ENDS

.subckt control_logic_delay_chain4 din dout vdd vss
Xinv0 din tmp0 vdd vss control_logic_inv
Xinv1 tmp0 tmp1 vdd vss control_logic_inv
Xinv2 tmp1 tmp2 vdd vss control_logic_inv
Xinv3 tmp2 dout vdd vss control_logic_inv
.ends

.subckt control_logic_delay_chain7 din dout vdd vss
Xinv0 din tmp0 vdd vss control_logic_inv
Xinv1 tmp0 tmp1 vdd vss control_logic_inv
Xinv2 tmp1 tmp2 vdd vss control_logic_inv
Xinv3 tmp2 tmp3 vdd vss control_logic_inv
Xinv4 tmp3 tmp4 vdd vss control_logic_inv
Xinv5 tmp4 tmp5 vdd vss control_logic_inv
Xinv6 tmp5 dout vdd vss control_logic_inv
.ends

.subckt control_logic_delay_chain8 din dout vdd vss
Xinv0 din tmp0 vdd vss control_logic_inv
Xinv1 tmp0 tmp1 vdd vss control_logic_inv
Xinv2 tmp1 tmp2 vdd vss control_logic_inv
Xinv3 tmp2 tmp3 vdd vss control_logic_inv
Xinv4 tmp3 tmp4 vdd vss control_logic_inv
Xinv5 tmp4 tmp5 vdd vss control_logic_inv
Xinv6 tmp5 tmp6 vdd vss control_logic_inv
Xinv7 tmp6 dout vdd vss control_logic_inv
.ends

.subckt control_logic_delay_chain16 din dout vdd vss
Xinv0 din tmp0 vdd vss control_logic_inv
Xinv1 tmp0 tmp1 vdd vss control_logic_inv
Xinv2 tmp1 tmp2 vdd vss control_logic_inv
Xinv3 tmp2 tmp3 vdd vss control_logic_inv
Xinv4 tmp3 tmp4 vdd vss control_logic_inv
Xinv5 tmp4 tmp5 vdd vss control_logic_inv
Xinv6 tmp5 tmp6 vdd vss control_logic_inv
Xinv7 tmp6 tmp7 vdd vss control_logic_inv
Xinv8 tmp7 tmp8 vdd vss control_logic_inv
Xinv9 tmp8 tmp9 vdd vss control_logic_inv
Xinv10 tmp9 tmp10 vdd vss control_logic_inv
Xinv11 tmp10 tmp11 vdd vss control_logic_inv
Xinv12 tmp11 tmp12 vdd vss control_logic_inv
Xinv13 tmp12 tmp13 vdd vss control_logic_inv
Xinv14 tmp13 tmp14 vdd vss control_logic_inv
Xinv15 tmp14 dout vdd vss control_logic_inv
.ends

.subckt control_logic_mux2 A0 A1 S X VPWR VGND
X0 a_27_368# A0 a_116_368# VPWR sky130_fd_pr__pfet_01v8 w=1 l=0.15
X1 a_27_368# S VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 X a_116_368# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_116_368# X VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_459_48# a_38_74# VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_459_48# S VPWR VPWR sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 X a_116_368# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=0.15
X7 a_270_74# S VGND VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_459_48# S VGND VGND sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 a_116_368# A1 a_206_368# VPWR sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR a_116_368# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=0.15
X11 VPWR a_459_48# a_206_368# VPWR sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_38_74# A0 a_116_368# VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_116_368# A1 a_270_74# VGND sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends

.subckt control_logic_bufbuf_16 A X VPWR VGND
X0 a_27_368# A VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_203_74# a_27_368# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND a_203_74# a_588_74# VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_203_74# a_588_74# VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_203_74# a_588_74# VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_588_74# a_203_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_588_74# a_203_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_588_74# a_203_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_588_74# a_203_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_588_74# a_203_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR a_203_74# a_588_74# VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_27_368# A VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_588_74# a_203_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VPWR a_27_368# a_203_74# VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR a_27_368# a_203_74# VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X35 VPWR a_203_74# a_588_74# VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X36 a_203_74# a_27_368# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X41 VPWR a_588_74# X VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X42 VPWR a_203_74# a_588_74# VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X43 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X44 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X45 VGND a_27_368# a_203_74# VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X46 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X47 VGND a_27_368# a_203_74# VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X48 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X49 VGND a_588_74# X VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X50 X a_588_74# VPWR VPWR sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X51 X a_588_74# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

.subckt control_logic_edge_detector din dout vdd vss 
xdelay_chain 
+ din delayed vdd vss 
+ control_logic_delay_chain7 

xand 
+ din delayed dout vdd vss 
+ control_logic_and2
.ends

.subckt sramgen_control_logic_replica_v2 clk we rbl dummy_bl pc_b wl_en0 wl_en write_driver_en sense_en vdd vss
* INPUT: clk we
* INOUT: rbl dummy_bl vdd vss
* OUTPUT: pc_b wl_en0 wl_en write_driver_en sense_en
Xinv_clk clk clk_b vdd vss control_logic_inv
Xinv_clk_b clk_b clk_buf vdd vss control_logic_inv
Xclk_pulse clk_buf clkp vdd vss control_logic_edge_detector
Xdecoder_replica clkp wl_en_set vdd vss control_logic_delay_chain8
Xinv_we we we_b vdd vss control_logic_inv

* Turn on wordlines at start of cycle
* Turn them off when replica bitline drops low enough
* to flip an inverter.
Xinv_rbl rbl rbl_b vdd vss control_logic_inv
Xpc_read_set_buf rbl_b pc_read_set vdd vss control_logic_delay_chain4
Xand_sense_en we_b rbl_b sense_en_set vdd vss control_logic_and2

Xwl_ctl wl_en_set wl_en_rst wl_en0 wl_en0_b vdd vss control_logic_sr_latch
Xsae_ctl sense_en_set clkp sense_en0 sense_en_b vdd vss control_logic_sr_latch
Xpc_ctl pc_set clkp pc pc_b0 vdd vss control_logic_sr_latch
Xwr_drv_ctl wr_drv_set wl_en_write_rst write_driver_en0 write_driver_en_b vdd vss control_logic_sr_latch

Xmux_wl_en_rst rbl_b wl_en_write_rst we wl_en_rst vdd vss control_logic_mux2
Xmux_pc_set pc_read_set pc_write_set we pc_set vdd vss control_logic_mux2
Xsae_set we_b rbl_b sae_set vdd vss control_logic_and2

Xwr_drv_set clkp we wr_drv_set vdd vss control_logic_and2
Xinv_dummy_bl dummy_bl dummy_bl_b vdd vss control_logic_inv
Xwl_en_write_rst_buf dummy_bl_b wl_en_write_rst vdd vss control_logic_delay_chain4
Xpc_write_set_buf wl_en_write_rst pc_write_set vdd vss control_logic_delay_chain4

Xwl_en_buf wl_en0 wl_en vdd vss control_logic_bufbuf_16
Xsae_buf sense_en0 sense_en vdd vss control_logic_bufbuf_16
Xpc_b_buf pc_b0 pc_b vdd vss control_logic_bufbuf_16
Xwr_drv_buf write_driver_en0 write_driver_en vdd vss control_logic_bufbuf_16

Xdummy_bl_pulldown dummy_bl write_driver_en0 vss vss sky130_fd_pr__nfet_01v8 w=0.800 l=0.150
.ends

