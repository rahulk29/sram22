magic
tech sky130A
magscale 1 2
timestamp 1623956458
<< nwell >>
rect 1558 428 1937 429
rect 886 -106 1937 428
<< pwell >>
rect 366 289 449 343
<< nmos >>
rect 92 159 240 189
rect 600 204 748 234
rect 600 132 748 162
rect 92 87 240 117
<< pmos >>
rect 1056 187 1280 217
rect 1522 186 1746 216
rect 1056 87 1280 117
rect 1522 87 1746 117
<< ndiff >>
rect 600 281 748 289
rect 92 238 240 246
rect 92 204 149 238
rect 183 204 240 238
rect 92 189 240 204
rect 600 247 663 281
rect 697 247 748 281
rect 600 234 748 247
rect 92 117 240 159
rect 600 162 748 204
rect 600 121 748 132
rect 92 71 240 87
rect 92 37 146 71
rect 180 37 240 71
rect 92 27 240 37
rect 600 87 661 121
rect 695 87 748 121
rect 600 79 748 87
<< pdiff >>
rect 1056 269 1280 277
rect 1056 235 1151 269
rect 1185 235 1280 269
rect 1056 217 1280 235
rect 1522 266 1746 277
rect 1522 232 1617 266
rect 1651 232 1746 266
rect 1522 216 1746 232
rect 1056 169 1280 187
rect 1056 135 1151 169
rect 1185 135 1280 169
rect 1056 117 1280 135
rect 1522 169 1746 186
rect 1522 135 1617 169
rect 1651 135 1746 169
rect 1522 117 1746 135
rect 1056 76 1280 87
rect 1056 42 1151 76
rect 1185 42 1280 76
rect 1056 27 1280 42
rect 1522 76 1746 87
rect 1522 42 1617 76
rect 1651 42 1746 76
rect 1522 27 1746 42
<< ndiffc >>
rect 149 204 183 238
rect 663 247 697 281
rect 146 37 180 71
rect 661 87 695 121
<< pdiffc >>
rect 1151 235 1185 269
rect 1617 232 1651 266
rect 1151 135 1185 169
rect 1617 135 1651 169
rect 1151 42 1185 76
rect 1617 42 1651 76
<< psubdiff >>
rect 366 333 449 343
rect 366 299 390 333
rect 424 299 449 333
rect 366 289 449 299
<< nsubdiff >>
rect 1807 230 1833 264
rect 1867 230 1900 264
<< psubdiffcont >>
rect 390 299 424 333
<< nsubdiffcont >>
rect 1833 230 1867 264
<< poly >>
rect 0 285 68 295
rect 0 251 17 285
rect 51 251 68 285
rect 0 189 68 251
rect 518 254 572 270
rect 278 222 334 238
rect 278 190 289 222
rect 273 189 289 190
rect 0 159 92 189
rect 240 188 289 189
rect 323 188 334 222
rect 518 220 528 254
rect 562 234 572 254
rect 803 254 858 270
rect 803 234 814 254
rect 562 220 600 234
rect 518 204 600 220
rect 748 220 814 234
rect 848 220 858 254
rect 748 204 858 220
rect 1400 276 1454 292
rect 1400 242 1410 276
rect 1444 242 1454 276
rect 240 159 334 188
rect 408 178 476 194
rect 408 144 418 178
rect 452 162 476 178
rect 905 187 1056 217
rect 1280 187 1306 217
rect 1400 210 1454 242
rect 905 162 935 187
rect 452 144 600 162
rect 408 132 600 144
rect 748 132 935 162
rect 408 128 476 132
rect 0 87 92 117
rect 240 87 359 117
rect 0 70 66 87
rect 0 36 16 70
rect 50 36 66 70
rect 0 26 66 36
rect 329 64 359 87
rect 1412 117 1442 210
rect 1496 186 1522 216
rect 1746 186 1867 216
rect 1813 181 1867 186
rect 1813 147 1823 181
rect 1857 147 1867 181
rect 1813 131 1867 147
rect 982 90 1056 117
rect 856 87 1056 90
rect 1280 87 1306 117
rect 1412 87 1522 117
rect 1746 87 1773 117
rect 856 64 1016 87
rect 329 60 1016 64
rect 329 34 886 60
<< polycont >>
rect 17 251 51 285
rect 289 188 323 222
rect 528 220 562 254
rect 814 220 848 254
rect 1410 242 1444 276
rect 418 144 452 178
rect 16 36 50 70
rect 1823 147 1857 181
<< locali >>
rect 135 333 457 343
rect 135 299 390 333
rect 424 299 457 333
rect 135 291 457 299
rect 0 251 17 285
rect 51 251 68 285
rect 135 241 182 291
rect 340 281 457 291
rect 612 281 744 284
rect 103 238 230 241
rect 0 214 66 217
rect 0 180 20 214
rect 54 180 66 214
rect 103 204 142 238
rect 183 204 230 238
rect 103 202 230 204
rect 273 222 341 224
rect 0 176 66 180
rect 273 177 289 222
rect 323 177 341 222
rect 512 220 528 254
rect 562 220 578 254
rect 612 247 663 281
rect 697 247 744 281
rect 1394 276 1479 278
rect 983 269 1159 270
rect 612 245 744 247
rect 798 254 883 256
rect 798 209 814 254
rect 848 214 883 254
rect 983 236 1151 269
rect 848 209 866 214
rect 798 197 866 209
rect 273 176 341 177
rect 402 178 470 196
rect 402 144 418 178
rect 452 144 470 178
rect 402 142 470 144
rect 0 108 470 142
rect 983 122 1017 236
rect 1134 235 1151 236
rect 1185 235 1202 269
rect 1394 231 1410 276
rect 1444 236 1479 276
rect 1444 231 1462 236
rect 1601 232 1617 266
rect 1651 232 1735 266
rect 1394 219 1462 231
rect 1134 135 1151 169
rect 1185 135 1617 169
rect 1651 135 1667 169
rect 614 121 1017 122
rect 614 87 661 121
rect 695 88 1017 121
rect 695 87 748 88
rect 983 76 1017 88
rect 1701 76 1735 232
rect 1807 230 1832 264
rect 1867 230 1900 264
rect 1807 181 1875 183
rect 1807 136 1823 181
rect 1857 136 1875 181
rect 1807 124 1875 136
rect 103 71 304 74
rect 0 36 16 70
rect 50 36 66 70
rect 103 37 146 71
rect 180 37 262 71
rect 296 37 304 71
rect 983 42 1151 76
rect 1185 42 1617 76
rect 1651 42 1828 76
rect 103 35 304 37
<< viali >>
rect 20 180 54 214
rect 142 204 149 238
rect 149 204 176 238
rect 289 188 323 211
rect 289 177 323 188
rect 528 220 562 254
rect 663 247 697 281
rect 814 220 848 243
rect 814 209 848 220
rect 418 144 452 178
rect 1410 242 1444 265
rect 1410 231 1444 242
rect 1151 135 1185 169
rect 1617 135 1651 169
rect 1832 230 1833 264
rect 1833 230 1866 264
rect 1823 147 1857 170
rect 1823 136 1857 147
rect 262 37 296 71
<< metal1 >>
rect 135 238 182 320
rect 656 281 706 293
rect 1 220 68 224
rect 1 168 7 220
rect 59 168 68 220
rect 135 204 142 238
rect 176 204 182 238
rect 514 264 578 270
rect 135 191 182 204
rect 273 219 341 224
rect 1 162 68 168
rect 273 167 281 219
rect 333 212 341 219
rect 514 212 520 264
rect 572 212 578 264
rect 656 247 663 281
rect 697 247 706 281
rect 656 240 706 247
rect 798 244 866 256
rect 798 243 867 244
rect 798 240 814 243
rect 848 240 867 243
rect 333 167 342 212
rect 514 206 578 212
rect 273 160 342 167
rect 406 178 470 196
rect 406 144 418 178
rect 452 144 470 178
rect 406 132 470 144
rect 243 71 311 83
rect 243 37 262 71
rect 296 57 311 71
rect 663 57 697 240
rect 798 188 806 240
rect 858 188 867 240
rect 798 181 867 188
rect 296 37 697 57
rect 243 29 697 37
rect 1144 169 1192 322
rect 1610 280 1658 321
rect 1394 266 1462 278
rect 1394 265 1463 266
rect 1394 262 1410 265
rect 1444 262 1463 265
rect 1394 210 1402 262
rect 1454 210 1463 262
rect 1394 203 1463 210
rect 1610 264 1904 280
rect 1610 232 1832 264
rect 1144 135 1151 169
rect 1185 135 1192 169
rect 1144 -32 1192 135
rect 1610 169 1658 232
rect 1825 230 1832 232
rect 1866 232 1904 264
rect 1866 230 1873 232
rect 1825 214 1873 230
rect 1610 135 1617 169
rect 1651 135 1658 169
rect 1610 -32 1658 135
rect 1807 170 1875 183
rect 1807 167 1823 170
rect 1857 167 1875 170
rect 1807 115 1815 167
rect 1867 115 1875 167
rect 1807 108 1875 115
<< via1 >>
rect 7 214 59 220
rect 7 180 20 214
rect 20 180 54 214
rect 54 180 59 214
rect 7 168 59 180
rect 281 211 333 219
rect 520 254 572 264
rect 520 220 528 254
rect 528 220 562 254
rect 562 220 572 254
rect 520 212 572 220
rect 281 177 289 211
rect 289 177 323 211
rect 323 177 333 211
rect 281 167 333 177
rect 806 209 814 240
rect 814 209 848 240
rect 848 209 858 240
rect 806 188 858 209
rect 1402 231 1410 262
rect 1410 231 1444 262
rect 1444 231 1454 262
rect 1402 210 1454 231
rect 1815 136 1823 167
rect 1823 136 1857 167
rect 1857 136 1867 167
rect 1815 115 1867 136
<< metal2 >>
rect 217 264 578 280
rect 217 252 520 264
rect 1 220 68 224
rect 1 168 7 220
rect 59 190 68 220
rect 217 190 245 252
rect 59 168 245 190
rect 1 162 245 168
rect 273 219 341 224
rect 273 167 281 219
rect 333 196 341 219
rect 514 212 520 252
rect 572 212 578 264
rect 954 262 1481 264
rect 954 242 1402 262
rect 514 206 578 212
rect 798 240 1402 242
rect 333 167 340 196
rect 798 188 806 240
rect 858 236 1402 240
rect 858 214 982 236
rect 858 188 867 214
rect 1394 210 1402 236
rect 1454 236 1481 262
rect 1454 210 1463 236
rect 1394 203 1463 210
rect 798 181 867 188
rect 273 159 340 167
rect 308 113 340 159
rect 1794 167 1875 184
rect 1794 115 1815 167
rect 1867 115 1875 167
rect 1794 113 1875 115
rect 308 108 1875 113
rect 308 85 1822 108
<< labels >>
rlabel metal1 s 135 185 182 320 4 GND
rlabel metal1 s 1610 -32 1658 231 4 VDD
rlabel metal1 s 158 252 158 252 4 gnd
rlabel polycont 34 268 34 268 1 A
rlabel locali 0 196 0 196 3 B
rlabel locali 1 126 1 126 3 C
rlabel polycont 33 53 33 53 1 D
rlabel metal1 s 1634 126 1634 126 4 vdd
rlabel metal1 s 1634 100 1634 100 4 vdd
rlabel locali 1798 60 1798 60 1 Z
rlabel metal1 s 1168 151 1168 151 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1937 316
<< end >>
